magic
tech gf180mcuD
magscale 1 5
timestamp 1701983776
<< obsm1 >>
rect 672 855 88648 89406
<< metal2 >>
rect 10976 0 11032 400
rect 11200 0 11256 400
rect 11424 0 11480 400
rect 11648 0 11704 400
rect 11872 0 11928 400
rect 12096 0 12152 400
rect 12320 0 12376 400
rect 12544 0 12600 400
rect 12768 0 12824 400
rect 12992 0 13048 400
rect 13216 0 13272 400
rect 13440 0 13496 400
rect 13664 0 13720 400
rect 13888 0 13944 400
rect 14112 0 14168 400
rect 14336 0 14392 400
rect 14560 0 14616 400
rect 14784 0 14840 400
rect 15008 0 15064 400
rect 15232 0 15288 400
rect 15456 0 15512 400
rect 15680 0 15736 400
rect 15904 0 15960 400
rect 16128 0 16184 400
rect 16352 0 16408 400
rect 16576 0 16632 400
rect 16800 0 16856 400
rect 17024 0 17080 400
rect 17248 0 17304 400
rect 17472 0 17528 400
rect 17696 0 17752 400
rect 17920 0 17976 400
rect 18144 0 18200 400
rect 18368 0 18424 400
rect 18592 0 18648 400
rect 18816 0 18872 400
rect 19040 0 19096 400
rect 19264 0 19320 400
rect 19488 0 19544 400
rect 19712 0 19768 400
rect 19936 0 19992 400
rect 20160 0 20216 400
rect 20384 0 20440 400
rect 20608 0 20664 400
rect 20832 0 20888 400
rect 21056 0 21112 400
rect 21280 0 21336 400
rect 21504 0 21560 400
rect 21728 0 21784 400
rect 21952 0 22008 400
rect 22176 0 22232 400
rect 22400 0 22456 400
rect 22624 0 22680 400
rect 22848 0 22904 400
rect 23072 0 23128 400
rect 23296 0 23352 400
rect 23520 0 23576 400
rect 23744 0 23800 400
rect 23968 0 24024 400
rect 24192 0 24248 400
rect 24416 0 24472 400
rect 24640 0 24696 400
rect 24864 0 24920 400
rect 25088 0 25144 400
rect 25312 0 25368 400
rect 25536 0 25592 400
rect 25760 0 25816 400
rect 25984 0 26040 400
rect 26208 0 26264 400
rect 26432 0 26488 400
rect 26656 0 26712 400
rect 26880 0 26936 400
rect 27104 0 27160 400
rect 27328 0 27384 400
rect 27552 0 27608 400
rect 27776 0 27832 400
rect 28000 0 28056 400
rect 28224 0 28280 400
rect 28448 0 28504 400
rect 28672 0 28728 400
rect 28896 0 28952 400
rect 29120 0 29176 400
rect 29344 0 29400 400
rect 29568 0 29624 400
rect 29792 0 29848 400
rect 30016 0 30072 400
rect 30240 0 30296 400
rect 30464 0 30520 400
rect 30688 0 30744 400
rect 30912 0 30968 400
rect 31136 0 31192 400
rect 31360 0 31416 400
rect 31584 0 31640 400
rect 31808 0 31864 400
rect 32032 0 32088 400
rect 32256 0 32312 400
rect 32480 0 32536 400
rect 32704 0 32760 400
rect 32928 0 32984 400
rect 33152 0 33208 400
rect 33376 0 33432 400
rect 33600 0 33656 400
rect 33824 0 33880 400
rect 34048 0 34104 400
rect 34272 0 34328 400
rect 34496 0 34552 400
rect 34720 0 34776 400
rect 34944 0 35000 400
rect 35168 0 35224 400
rect 35392 0 35448 400
rect 35616 0 35672 400
rect 35840 0 35896 400
rect 36064 0 36120 400
rect 36288 0 36344 400
rect 36512 0 36568 400
rect 36736 0 36792 400
rect 36960 0 37016 400
rect 37184 0 37240 400
rect 37408 0 37464 400
rect 37632 0 37688 400
rect 37856 0 37912 400
rect 38080 0 38136 400
rect 38304 0 38360 400
rect 38528 0 38584 400
rect 38752 0 38808 400
rect 38976 0 39032 400
rect 39200 0 39256 400
rect 39424 0 39480 400
rect 39648 0 39704 400
rect 39872 0 39928 400
rect 40096 0 40152 400
rect 40320 0 40376 400
rect 40544 0 40600 400
rect 40768 0 40824 400
rect 40992 0 41048 400
rect 41216 0 41272 400
rect 41440 0 41496 400
rect 41664 0 41720 400
rect 41888 0 41944 400
rect 42112 0 42168 400
rect 42336 0 42392 400
rect 42560 0 42616 400
rect 42784 0 42840 400
rect 43008 0 43064 400
rect 43232 0 43288 400
rect 43456 0 43512 400
rect 43680 0 43736 400
rect 43904 0 43960 400
rect 44128 0 44184 400
rect 44352 0 44408 400
rect 44576 0 44632 400
rect 44800 0 44856 400
rect 45024 0 45080 400
rect 45248 0 45304 400
rect 45472 0 45528 400
rect 45696 0 45752 400
rect 45920 0 45976 400
rect 46144 0 46200 400
rect 46368 0 46424 400
rect 46592 0 46648 400
rect 46816 0 46872 400
rect 47040 0 47096 400
rect 47264 0 47320 400
rect 47488 0 47544 400
rect 47712 0 47768 400
rect 47936 0 47992 400
rect 48160 0 48216 400
rect 48384 0 48440 400
rect 48608 0 48664 400
rect 48832 0 48888 400
rect 49056 0 49112 400
rect 49280 0 49336 400
rect 49504 0 49560 400
rect 49728 0 49784 400
rect 49952 0 50008 400
rect 50176 0 50232 400
rect 50400 0 50456 400
rect 50624 0 50680 400
rect 50848 0 50904 400
rect 51072 0 51128 400
rect 51296 0 51352 400
rect 51520 0 51576 400
rect 51744 0 51800 400
rect 51968 0 52024 400
rect 52192 0 52248 400
rect 52416 0 52472 400
rect 52640 0 52696 400
rect 52864 0 52920 400
rect 53088 0 53144 400
rect 53312 0 53368 400
rect 53536 0 53592 400
rect 53760 0 53816 400
rect 53984 0 54040 400
rect 54208 0 54264 400
rect 54432 0 54488 400
rect 54656 0 54712 400
rect 54880 0 54936 400
rect 55104 0 55160 400
rect 55328 0 55384 400
rect 55552 0 55608 400
rect 55776 0 55832 400
rect 56000 0 56056 400
rect 56224 0 56280 400
rect 56448 0 56504 400
rect 56672 0 56728 400
rect 56896 0 56952 400
rect 57120 0 57176 400
rect 57344 0 57400 400
rect 57568 0 57624 400
rect 57792 0 57848 400
rect 58016 0 58072 400
rect 58240 0 58296 400
rect 58464 0 58520 400
rect 58688 0 58744 400
rect 58912 0 58968 400
rect 59136 0 59192 400
rect 59360 0 59416 400
rect 59584 0 59640 400
rect 59808 0 59864 400
rect 60032 0 60088 400
rect 60256 0 60312 400
rect 60480 0 60536 400
rect 60704 0 60760 400
rect 60928 0 60984 400
rect 61152 0 61208 400
rect 61376 0 61432 400
rect 61600 0 61656 400
rect 61824 0 61880 400
rect 62048 0 62104 400
rect 62272 0 62328 400
rect 62496 0 62552 400
rect 62720 0 62776 400
rect 62944 0 63000 400
rect 63168 0 63224 400
rect 63392 0 63448 400
rect 63616 0 63672 400
rect 63840 0 63896 400
rect 64064 0 64120 400
rect 64288 0 64344 400
rect 64512 0 64568 400
rect 64736 0 64792 400
rect 64960 0 65016 400
rect 65184 0 65240 400
rect 65408 0 65464 400
rect 65632 0 65688 400
rect 65856 0 65912 400
rect 66080 0 66136 400
rect 66304 0 66360 400
rect 66528 0 66584 400
rect 66752 0 66808 400
rect 66976 0 67032 400
rect 67200 0 67256 400
rect 67424 0 67480 400
rect 67648 0 67704 400
rect 67872 0 67928 400
rect 68096 0 68152 400
rect 68320 0 68376 400
rect 68544 0 68600 400
rect 68768 0 68824 400
rect 68992 0 69048 400
rect 69216 0 69272 400
rect 69440 0 69496 400
rect 69664 0 69720 400
rect 69888 0 69944 400
rect 70112 0 70168 400
rect 70336 0 70392 400
rect 70560 0 70616 400
rect 70784 0 70840 400
rect 71008 0 71064 400
rect 71232 0 71288 400
rect 71456 0 71512 400
rect 71680 0 71736 400
rect 71904 0 71960 400
rect 72128 0 72184 400
rect 72352 0 72408 400
rect 72576 0 72632 400
rect 72800 0 72856 400
rect 73024 0 73080 400
rect 73248 0 73304 400
rect 73472 0 73528 400
rect 73696 0 73752 400
rect 73920 0 73976 400
rect 74144 0 74200 400
rect 74368 0 74424 400
rect 74592 0 74648 400
rect 74816 0 74872 400
rect 75040 0 75096 400
rect 75264 0 75320 400
rect 75488 0 75544 400
rect 75712 0 75768 400
rect 75936 0 75992 400
rect 76160 0 76216 400
rect 76384 0 76440 400
rect 76608 0 76664 400
rect 76832 0 76888 400
rect 77056 0 77112 400
rect 77280 0 77336 400
rect 77504 0 77560 400
rect 77728 0 77784 400
rect 77952 0 78008 400
rect 78176 0 78232 400
<< obsm2 >>
rect 574 430 88858 89395
rect 574 400 10946 430
rect 11062 400 11170 430
rect 11286 400 11394 430
rect 11510 400 11618 430
rect 11734 400 11842 430
rect 11958 400 12066 430
rect 12182 400 12290 430
rect 12406 400 12514 430
rect 12630 400 12738 430
rect 12854 400 12962 430
rect 13078 400 13186 430
rect 13302 400 13410 430
rect 13526 400 13634 430
rect 13750 400 13858 430
rect 13974 400 14082 430
rect 14198 400 14306 430
rect 14422 400 14530 430
rect 14646 400 14754 430
rect 14870 400 14978 430
rect 15094 400 15202 430
rect 15318 400 15426 430
rect 15542 400 15650 430
rect 15766 400 15874 430
rect 15990 400 16098 430
rect 16214 400 16322 430
rect 16438 400 16546 430
rect 16662 400 16770 430
rect 16886 400 16994 430
rect 17110 400 17218 430
rect 17334 400 17442 430
rect 17558 400 17666 430
rect 17782 400 17890 430
rect 18006 400 18114 430
rect 18230 400 18338 430
rect 18454 400 18562 430
rect 18678 400 18786 430
rect 18902 400 19010 430
rect 19126 400 19234 430
rect 19350 400 19458 430
rect 19574 400 19682 430
rect 19798 400 19906 430
rect 20022 400 20130 430
rect 20246 400 20354 430
rect 20470 400 20578 430
rect 20694 400 20802 430
rect 20918 400 21026 430
rect 21142 400 21250 430
rect 21366 400 21474 430
rect 21590 400 21698 430
rect 21814 400 21922 430
rect 22038 400 22146 430
rect 22262 400 22370 430
rect 22486 400 22594 430
rect 22710 400 22818 430
rect 22934 400 23042 430
rect 23158 400 23266 430
rect 23382 400 23490 430
rect 23606 400 23714 430
rect 23830 400 23938 430
rect 24054 400 24162 430
rect 24278 400 24386 430
rect 24502 400 24610 430
rect 24726 400 24834 430
rect 24950 400 25058 430
rect 25174 400 25282 430
rect 25398 400 25506 430
rect 25622 400 25730 430
rect 25846 400 25954 430
rect 26070 400 26178 430
rect 26294 400 26402 430
rect 26518 400 26626 430
rect 26742 400 26850 430
rect 26966 400 27074 430
rect 27190 400 27298 430
rect 27414 400 27522 430
rect 27638 400 27746 430
rect 27862 400 27970 430
rect 28086 400 28194 430
rect 28310 400 28418 430
rect 28534 400 28642 430
rect 28758 400 28866 430
rect 28982 400 29090 430
rect 29206 400 29314 430
rect 29430 400 29538 430
rect 29654 400 29762 430
rect 29878 400 29986 430
rect 30102 400 30210 430
rect 30326 400 30434 430
rect 30550 400 30658 430
rect 30774 400 30882 430
rect 30998 400 31106 430
rect 31222 400 31330 430
rect 31446 400 31554 430
rect 31670 400 31778 430
rect 31894 400 32002 430
rect 32118 400 32226 430
rect 32342 400 32450 430
rect 32566 400 32674 430
rect 32790 400 32898 430
rect 33014 400 33122 430
rect 33238 400 33346 430
rect 33462 400 33570 430
rect 33686 400 33794 430
rect 33910 400 34018 430
rect 34134 400 34242 430
rect 34358 400 34466 430
rect 34582 400 34690 430
rect 34806 400 34914 430
rect 35030 400 35138 430
rect 35254 400 35362 430
rect 35478 400 35586 430
rect 35702 400 35810 430
rect 35926 400 36034 430
rect 36150 400 36258 430
rect 36374 400 36482 430
rect 36598 400 36706 430
rect 36822 400 36930 430
rect 37046 400 37154 430
rect 37270 400 37378 430
rect 37494 400 37602 430
rect 37718 400 37826 430
rect 37942 400 38050 430
rect 38166 400 38274 430
rect 38390 400 38498 430
rect 38614 400 38722 430
rect 38838 400 38946 430
rect 39062 400 39170 430
rect 39286 400 39394 430
rect 39510 400 39618 430
rect 39734 400 39842 430
rect 39958 400 40066 430
rect 40182 400 40290 430
rect 40406 400 40514 430
rect 40630 400 40738 430
rect 40854 400 40962 430
rect 41078 400 41186 430
rect 41302 400 41410 430
rect 41526 400 41634 430
rect 41750 400 41858 430
rect 41974 400 42082 430
rect 42198 400 42306 430
rect 42422 400 42530 430
rect 42646 400 42754 430
rect 42870 400 42978 430
rect 43094 400 43202 430
rect 43318 400 43426 430
rect 43542 400 43650 430
rect 43766 400 43874 430
rect 43990 400 44098 430
rect 44214 400 44322 430
rect 44438 400 44546 430
rect 44662 400 44770 430
rect 44886 400 44994 430
rect 45110 400 45218 430
rect 45334 400 45442 430
rect 45558 400 45666 430
rect 45782 400 45890 430
rect 46006 400 46114 430
rect 46230 400 46338 430
rect 46454 400 46562 430
rect 46678 400 46786 430
rect 46902 400 47010 430
rect 47126 400 47234 430
rect 47350 400 47458 430
rect 47574 400 47682 430
rect 47798 400 47906 430
rect 48022 400 48130 430
rect 48246 400 48354 430
rect 48470 400 48578 430
rect 48694 400 48802 430
rect 48918 400 49026 430
rect 49142 400 49250 430
rect 49366 400 49474 430
rect 49590 400 49698 430
rect 49814 400 49922 430
rect 50038 400 50146 430
rect 50262 400 50370 430
rect 50486 400 50594 430
rect 50710 400 50818 430
rect 50934 400 51042 430
rect 51158 400 51266 430
rect 51382 400 51490 430
rect 51606 400 51714 430
rect 51830 400 51938 430
rect 52054 400 52162 430
rect 52278 400 52386 430
rect 52502 400 52610 430
rect 52726 400 52834 430
rect 52950 400 53058 430
rect 53174 400 53282 430
rect 53398 400 53506 430
rect 53622 400 53730 430
rect 53846 400 53954 430
rect 54070 400 54178 430
rect 54294 400 54402 430
rect 54518 400 54626 430
rect 54742 400 54850 430
rect 54966 400 55074 430
rect 55190 400 55298 430
rect 55414 400 55522 430
rect 55638 400 55746 430
rect 55862 400 55970 430
rect 56086 400 56194 430
rect 56310 400 56418 430
rect 56534 400 56642 430
rect 56758 400 56866 430
rect 56982 400 57090 430
rect 57206 400 57314 430
rect 57430 400 57538 430
rect 57654 400 57762 430
rect 57878 400 57986 430
rect 58102 400 58210 430
rect 58326 400 58434 430
rect 58550 400 58658 430
rect 58774 400 58882 430
rect 58998 400 59106 430
rect 59222 400 59330 430
rect 59446 400 59554 430
rect 59670 400 59778 430
rect 59894 400 60002 430
rect 60118 400 60226 430
rect 60342 400 60450 430
rect 60566 400 60674 430
rect 60790 400 60898 430
rect 61014 400 61122 430
rect 61238 400 61346 430
rect 61462 400 61570 430
rect 61686 400 61794 430
rect 61910 400 62018 430
rect 62134 400 62242 430
rect 62358 400 62466 430
rect 62582 400 62690 430
rect 62806 400 62914 430
rect 63030 400 63138 430
rect 63254 400 63362 430
rect 63478 400 63586 430
rect 63702 400 63810 430
rect 63926 400 64034 430
rect 64150 400 64258 430
rect 64374 400 64482 430
rect 64598 400 64706 430
rect 64822 400 64930 430
rect 65046 400 65154 430
rect 65270 400 65378 430
rect 65494 400 65602 430
rect 65718 400 65826 430
rect 65942 400 66050 430
rect 66166 400 66274 430
rect 66390 400 66498 430
rect 66614 400 66722 430
rect 66838 400 66946 430
rect 67062 400 67170 430
rect 67286 400 67394 430
rect 67510 400 67618 430
rect 67734 400 67842 430
rect 67958 400 68066 430
rect 68182 400 68290 430
rect 68406 400 68514 430
rect 68630 400 68738 430
rect 68854 400 68962 430
rect 69078 400 69186 430
rect 69302 400 69410 430
rect 69526 400 69634 430
rect 69750 400 69858 430
rect 69974 400 70082 430
rect 70198 400 70306 430
rect 70422 400 70530 430
rect 70646 400 70754 430
rect 70870 400 70978 430
rect 71094 400 71202 430
rect 71318 400 71426 430
rect 71542 400 71650 430
rect 71766 400 71874 430
rect 71990 400 72098 430
rect 72214 400 72322 430
rect 72438 400 72546 430
rect 72662 400 72770 430
rect 72886 400 72994 430
rect 73110 400 73218 430
rect 73334 400 73442 430
rect 73558 400 73666 430
rect 73782 400 73890 430
rect 74006 400 74114 430
rect 74230 400 74338 430
rect 74454 400 74562 430
rect 74678 400 74786 430
rect 74902 400 75010 430
rect 75126 400 75234 430
rect 75350 400 75458 430
rect 75574 400 75682 430
rect 75798 400 75906 430
rect 76022 400 76130 430
rect 76246 400 76354 430
rect 76470 400 76578 430
rect 76694 400 76802 430
rect 76918 400 77026 430
rect 77142 400 77250 430
rect 77366 400 77474 430
rect 77590 400 77698 430
rect 77814 400 77922 430
rect 78038 400 78146 430
rect 78262 400 88858 430
<< metal3 >>
rect 0 88032 400 88088
rect 88971 88032 89371 88088
rect 0 84336 400 84392
rect 88971 84336 89371 84392
rect 0 80640 400 80696
rect 88971 80640 89371 80696
rect 0 76944 400 77000
rect 88971 76944 89371 77000
rect 0 73248 400 73304
rect 88971 73248 89371 73304
rect 0 69552 400 69608
rect 88971 69552 89371 69608
rect 0 65856 400 65912
rect 88971 65856 89371 65912
rect 0 62160 400 62216
rect 88971 62160 89371 62216
rect 0 58464 400 58520
rect 88971 58464 89371 58520
rect 0 54768 400 54824
rect 88971 54768 89371 54824
rect 0 51072 400 51128
rect 88971 51072 89371 51128
rect 0 47376 400 47432
rect 88971 47376 89371 47432
rect 0 43680 400 43736
rect 88971 43680 89371 43736
rect 0 39984 400 40040
rect 88971 39984 89371 40040
rect 0 36288 400 36344
rect 88971 36288 89371 36344
rect 0 32592 400 32648
rect 88971 32592 89371 32648
rect 0 28896 400 28952
rect 88971 28896 89371 28952
rect 0 25200 400 25256
rect 88971 25200 89371 25256
rect 0 21504 400 21560
rect 88971 21504 89371 21560
rect 0 17808 400 17864
rect 88971 17808 89371 17864
rect 0 14112 400 14168
rect 88971 14112 89371 14168
rect 0 10416 400 10472
rect 88971 10416 89371 10472
rect 0 6720 400 6776
rect 88971 6720 89371 6776
rect 0 3024 400 3080
rect 88971 3024 89371 3080
<< obsm3 >>
rect 400 88118 88971 89390
rect 430 88002 88941 88118
rect 400 84422 88971 88002
rect 430 84306 88941 84422
rect 400 80726 88971 84306
rect 430 80610 88941 80726
rect 400 77030 88971 80610
rect 430 76914 88941 77030
rect 400 73334 88971 76914
rect 430 73218 88941 73334
rect 400 69638 88971 73218
rect 430 69522 88941 69638
rect 400 65942 88971 69522
rect 430 65826 88941 65942
rect 400 62246 88971 65826
rect 430 62130 88941 62246
rect 400 58550 88971 62130
rect 430 58434 88941 58550
rect 400 54854 88971 58434
rect 430 54738 88941 54854
rect 400 51158 88971 54738
rect 430 51042 88941 51158
rect 400 47462 88971 51042
rect 430 47346 88941 47462
rect 400 43766 88971 47346
rect 430 43650 88941 43766
rect 400 40070 88971 43650
rect 430 39954 88941 40070
rect 400 36374 88971 39954
rect 430 36258 88941 36374
rect 400 32678 88971 36258
rect 430 32562 88941 32678
rect 400 28982 88971 32562
rect 430 28866 88941 28982
rect 400 25286 88971 28866
rect 430 25170 88941 25286
rect 400 21590 88971 25170
rect 430 21474 88941 21590
rect 400 17894 88971 21474
rect 430 17778 88941 17894
rect 400 14198 88971 17778
rect 430 14082 88941 14198
rect 400 10502 88971 14082
rect 430 10386 88941 10502
rect 400 6806 88971 10386
rect 430 6690 88941 6806
rect 400 3110 88971 6690
rect 430 2994 88941 3110
rect 400 1358 88971 2994
<< metal4 >>
rect 2224 1538 2384 89406
rect 9904 1538 10064 89406
rect 17584 1538 17744 89406
rect 25264 1538 25424 89406
rect 32944 1538 33104 89406
rect 40624 1538 40784 89406
rect 48304 1538 48464 89406
rect 55984 1538 56144 89406
rect 63664 1538 63824 89406
rect 71344 1538 71504 89406
rect 79024 1538 79184 89406
rect 86704 1538 86864 89406
<< obsm4 >>
rect 1190 2529 2194 86511
rect 2414 2529 9874 86511
rect 10094 2529 17554 86511
rect 17774 2529 25234 86511
rect 25454 2529 32914 86511
rect 33134 2529 40594 86511
rect 40814 2529 48274 86511
rect 48494 2529 55954 86511
rect 56174 2529 63634 86511
rect 63854 2529 71314 86511
rect 71534 2529 78994 86511
rect 79214 2529 86674 86511
rect 86894 2529 88018 86511
<< labels >>
rlabel metal3 s 88971 3024 89371 3080 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 65856 400 65912 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 54768 400 54824 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 43680 400 43736 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 32592 400 32648 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 21504 400 21560 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 10416 400 10472 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 88971 14112 89371 14168 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 88971 25200 89371 25256 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 88971 36288 89371 36344 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 88971 47376 89371 47432 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 88971 58464 89371 58520 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 88971 69552 89371 69608 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 88971 80640 89371 80696 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 88032 400 88088 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 76944 400 77000 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 88971 10416 89371 10472 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 58464 400 58520 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 47376 400 47432 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 36288 400 36344 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 25200 400 25256 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 14112 400 14168 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 3024 400 3080 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 88971 21504 89371 21560 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 88971 32592 89371 32648 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 88971 43680 89371 43736 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 88971 54768 89371 54824 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 88971 65856 89371 65912 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 88971 76944 89371 77000 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 88971 88032 89371 88088 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 80640 400 80696 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 69552 400 69608 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 88971 6720 89371 6776 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 62160 400 62216 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 51072 400 51128 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 39984 400 40040 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 28896 400 28952 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 17808 400 17864 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 6720 400 6776 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 88971 17808 89371 17864 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 88971 28896 89371 28952 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 88971 39984 89371 40040 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 88971 51072 89371 51128 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 88971 62160 89371 62216 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 88971 73248 89371 73304 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 88971 84336 89371 84392 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 84336 400 84392 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 73248 400 73304 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 77728 0 77784 400 6 irq[0]
port 49 nsew signal output
rlabel metal2 s 77952 0 78008 400 6 irq[1]
port 50 nsew signal output
rlabel metal2 s 78176 0 78232 400 6 irq[2]
port 51 nsew signal output
rlabel metal2 s 34720 0 34776 400 6 la_data_in[0]
port 52 nsew signal input
rlabel metal2 s 41440 0 41496 400 6 la_data_in[10]
port 53 nsew signal input
rlabel metal2 s 42112 0 42168 400 6 la_data_in[11]
port 54 nsew signal input
rlabel metal2 s 42784 0 42840 400 6 la_data_in[12]
port 55 nsew signal input
rlabel metal2 s 43456 0 43512 400 6 la_data_in[13]
port 56 nsew signal input
rlabel metal2 s 44128 0 44184 400 6 la_data_in[14]
port 57 nsew signal input
rlabel metal2 s 44800 0 44856 400 6 la_data_in[15]
port 58 nsew signal input
rlabel metal2 s 45472 0 45528 400 6 la_data_in[16]
port 59 nsew signal input
rlabel metal2 s 46144 0 46200 400 6 la_data_in[17]
port 60 nsew signal input
rlabel metal2 s 46816 0 46872 400 6 la_data_in[18]
port 61 nsew signal input
rlabel metal2 s 47488 0 47544 400 6 la_data_in[19]
port 62 nsew signal input
rlabel metal2 s 35392 0 35448 400 6 la_data_in[1]
port 63 nsew signal input
rlabel metal2 s 48160 0 48216 400 6 la_data_in[20]
port 64 nsew signal input
rlabel metal2 s 48832 0 48888 400 6 la_data_in[21]
port 65 nsew signal input
rlabel metal2 s 49504 0 49560 400 6 la_data_in[22]
port 66 nsew signal input
rlabel metal2 s 50176 0 50232 400 6 la_data_in[23]
port 67 nsew signal input
rlabel metal2 s 50848 0 50904 400 6 la_data_in[24]
port 68 nsew signal input
rlabel metal2 s 51520 0 51576 400 6 la_data_in[25]
port 69 nsew signal input
rlabel metal2 s 52192 0 52248 400 6 la_data_in[26]
port 70 nsew signal input
rlabel metal2 s 52864 0 52920 400 6 la_data_in[27]
port 71 nsew signal input
rlabel metal2 s 53536 0 53592 400 6 la_data_in[28]
port 72 nsew signal input
rlabel metal2 s 54208 0 54264 400 6 la_data_in[29]
port 73 nsew signal input
rlabel metal2 s 36064 0 36120 400 6 la_data_in[2]
port 74 nsew signal input
rlabel metal2 s 54880 0 54936 400 6 la_data_in[30]
port 75 nsew signal input
rlabel metal2 s 55552 0 55608 400 6 la_data_in[31]
port 76 nsew signal input
rlabel metal2 s 56224 0 56280 400 6 la_data_in[32]
port 77 nsew signal input
rlabel metal2 s 56896 0 56952 400 6 la_data_in[33]
port 78 nsew signal input
rlabel metal2 s 57568 0 57624 400 6 la_data_in[34]
port 79 nsew signal input
rlabel metal2 s 58240 0 58296 400 6 la_data_in[35]
port 80 nsew signal input
rlabel metal2 s 58912 0 58968 400 6 la_data_in[36]
port 81 nsew signal input
rlabel metal2 s 59584 0 59640 400 6 la_data_in[37]
port 82 nsew signal input
rlabel metal2 s 60256 0 60312 400 6 la_data_in[38]
port 83 nsew signal input
rlabel metal2 s 60928 0 60984 400 6 la_data_in[39]
port 84 nsew signal input
rlabel metal2 s 36736 0 36792 400 6 la_data_in[3]
port 85 nsew signal input
rlabel metal2 s 61600 0 61656 400 6 la_data_in[40]
port 86 nsew signal input
rlabel metal2 s 62272 0 62328 400 6 la_data_in[41]
port 87 nsew signal input
rlabel metal2 s 62944 0 63000 400 6 la_data_in[42]
port 88 nsew signal input
rlabel metal2 s 63616 0 63672 400 6 la_data_in[43]
port 89 nsew signal input
rlabel metal2 s 64288 0 64344 400 6 la_data_in[44]
port 90 nsew signal input
rlabel metal2 s 64960 0 65016 400 6 la_data_in[45]
port 91 nsew signal input
rlabel metal2 s 65632 0 65688 400 6 la_data_in[46]
port 92 nsew signal input
rlabel metal2 s 66304 0 66360 400 6 la_data_in[47]
port 93 nsew signal input
rlabel metal2 s 66976 0 67032 400 6 la_data_in[48]
port 94 nsew signal input
rlabel metal2 s 67648 0 67704 400 6 la_data_in[49]
port 95 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 la_data_in[4]
port 96 nsew signal input
rlabel metal2 s 68320 0 68376 400 6 la_data_in[50]
port 97 nsew signal input
rlabel metal2 s 68992 0 69048 400 6 la_data_in[51]
port 98 nsew signal input
rlabel metal2 s 69664 0 69720 400 6 la_data_in[52]
port 99 nsew signal input
rlabel metal2 s 70336 0 70392 400 6 la_data_in[53]
port 100 nsew signal input
rlabel metal2 s 71008 0 71064 400 6 la_data_in[54]
port 101 nsew signal input
rlabel metal2 s 71680 0 71736 400 6 la_data_in[55]
port 102 nsew signal input
rlabel metal2 s 72352 0 72408 400 6 la_data_in[56]
port 103 nsew signal input
rlabel metal2 s 73024 0 73080 400 6 la_data_in[57]
port 104 nsew signal input
rlabel metal2 s 73696 0 73752 400 6 la_data_in[58]
port 105 nsew signal input
rlabel metal2 s 74368 0 74424 400 6 la_data_in[59]
port 106 nsew signal input
rlabel metal2 s 38080 0 38136 400 6 la_data_in[5]
port 107 nsew signal input
rlabel metal2 s 75040 0 75096 400 6 la_data_in[60]
port 108 nsew signal input
rlabel metal2 s 75712 0 75768 400 6 la_data_in[61]
port 109 nsew signal input
rlabel metal2 s 76384 0 76440 400 6 la_data_in[62]
port 110 nsew signal input
rlabel metal2 s 77056 0 77112 400 6 la_data_in[63]
port 111 nsew signal input
rlabel metal2 s 38752 0 38808 400 6 la_data_in[6]
port 112 nsew signal input
rlabel metal2 s 39424 0 39480 400 6 la_data_in[7]
port 113 nsew signal input
rlabel metal2 s 40096 0 40152 400 6 la_data_in[8]
port 114 nsew signal input
rlabel metal2 s 40768 0 40824 400 6 la_data_in[9]
port 115 nsew signal input
rlabel metal2 s 34944 0 35000 400 6 la_data_out[0]
port 116 nsew signal output
rlabel metal2 s 41664 0 41720 400 6 la_data_out[10]
port 117 nsew signal output
rlabel metal2 s 42336 0 42392 400 6 la_data_out[11]
port 118 nsew signal output
rlabel metal2 s 43008 0 43064 400 6 la_data_out[12]
port 119 nsew signal output
rlabel metal2 s 43680 0 43736 400 6 la_data_out[13]
port 120 nsew signal output
rlabel metal2 s 44352 0 44408 400 6 la_data_out[14]
port 121 nsew signal output
rlabel metal2 s 45024 0 45080 400 6 la_data_out[15]
port 122 nsew signal output
rlabel metal2 s 45696 0 45752 400 6 la_data_out[16]
port 123 nsew signal output
rlabel metal2 s 46368 0 46424 400 6 la_data_out[17]
port 124 nsew signal output
rlabel metal2 s 47040 0 47096 400 6 la_data_out[18]
port 125 nsew signal output
rlabel metal2 s 47712 0 47768 400 6 la_data_out[19]
port 126 nsew signal output
rlabel metal2 s 35616 0 35672 400 6 la_data_out[1]
port 127 nsew signal output
rlabel metal2 s 48384 0 48440 400 6 la_data_out[20]
port 128 nsew signal output
rlabel metal2 s 49056 0 49112 400 6 la_data_out[21]
port 129 nsew signal output
rlabel metal2 s 49728 0 49784 400 6 la_data_out[22]
port 130 nsew signal output
rlabel metal2 s 50400 0 50456 400 6 la_data_out[23]
port 131 nsew signal output
rlabel metal2 s 51072 0 51128 400 6 la_data_out[24]
port 132 nsew signal output
rlabel metal2 s 51744 0 51800 400 6 la_data_out[25]
port 133 nsew signal output
rlabel metal2 s 52416 0 52472 400 6 la_data_out[26]
port 134 nsew signal output
rlabel metal2 s 53088 0 53144 400 6 la_data_out[27]
port 135 nsew signal output
rlabel metal2 s 53760 0 53816 400 6 la_data_out[28]
port 136 nsew signal output
rlabel metal2 s 54432 0 54488 400 6 la_data_out[29]
port 137 nsew signal output
rlabel metal2 s 36288 0 36344 400 6 la_data_out[2]
port 138 nsew signal output
rlabel metal2 s 55104 0 55160 400 6 la_data_out[30]
port 139 nsew signal output
rlabel metal2 s 55776 0 55832 400 6 la_data_out[31]
port 140 nsew signal output
rlabel metal2 s 56448 0 56504 400 6 la_data_out[32]
port 141 nsew signal output
rlabel metal2 s 57120 0 57176 400 6 la_data_out[33]
port 142 nsew signal output
rlabel metal2 s 57792 0 57848 400 6 la_data_out[34]
port 143 nsew signal output
rlabel metal2 s 58464 0 58520 400 6 la_data_out[35]
port 144 nsew signal output
rlabel metal2 s 59136 0 59192 400 6 la_data_out[36]
port 145 nsew signal output
rlabel metal2 s 59808 0 59864 400 6 la_data_out[37]
port 146 nsew signal output
rlabel metal2 s 60480 0 60536 400 6 la_data_out[38]
port 147 nsew signal output
rlabel metal2 s 61152 0 61208 400 6 la_data_out[39]
port 148 nsew signal output
rlabel metal2 s 36960 0 37016 400 6 la_data_out[3]
port 149 nsew signal output
rlabel metal2 s 61824 0 61880 400 6 la_data_out[40]
port 150 nsew signal output
rlabel metal2 s 62496 0 62552 400 6 la_data_out[41]
port 151 nsew signal output
rlabel metal2 s 63168 0 63224 400 6 la_data_out[42]
port 152 nsew signal output
rlabel metal2 s 63840 0 63896 400 6 la_data_out[43]
port 153 nsew signal output
rlabel metal2 s 64512 0 64568 400 6 la_data_out[44]
port 154 nsew signal output
rlabel metal2 s 65184 0 65240 400 6 la_data_out[45]
port 155 nsew signal output
rlabel metal2 s 65856 0 65912 400 6 la_data_out[46]
port 156 nsew signal output
rlabel metal2 s 66528 0 66584 400 6 la_data_out[47]
port 157 nsew signal output
rlabel metal2 s 67200 0 67256 400 6 la_data_out[48]
port 158 nsew signal output
rlabel metal2 s 67872 0 67928 400 6 la_data_out[49]
port 159 nsew signal output
rlabel metal2 s 37632 0 37688 400 6 la_data_out[4]
port 160 nsew signal output
rlabel metal2 s 68544 0 68600 400 6 la_data_out[50]
port 161 nsew signal output
rlabel metal2 s 69216 0 69272 400 6 la_data_out[51]
port 162 nsew signal output
rlabel metal2 s 69888 0 69944 400 6 la_data_out[52]
port 163 nsew signal output
rlabel metal2 s 70560 0 70616 400 6 la_data_out[53]
port 164 nsew signal output
rlabel metal2 s 71232 0 71288 400 6 la_data_out[54]
port 165 nsew signal output
rlabel metal2 s 71904 0 71960 400 6 la_data_out[55]
port 166 nsew signal output
rlabel metal2 s 72576 0 72632 400 6 la_data_out[56]
port 167 nsew signal output
rlabel metal2 s 73248 0 73304 400 6 la_data_out[57]
port 168 nsew signal output
rlabel metal2 s 73920 0 73976 400 6 la_data_out[58]
port 169 nsew signal output
rlabel metal2 s 74592 0 74648 400 6 la_data_out[59]
port 170 nsew signal output
rlabel metal2 s 38304 0 38360 400 6 la_data_out[5]
port 171 nsew signal output
rlabel metal2 s 75264 0 75320 400 6 la_data_out[60]
port 172 nsew signal output
rlabel metal2 s 75936 0 75992 400 6 la_data_out[61]
port 173 nsew signal output
rlabel metal2 s 76608 0 76664 400 6 la_data_out[62]
port 174 nsew signal output
rlabel metal2 s 77280 0 77336 400 6 la_data_out[63]
port 175 nsew signal output
rlabel metal2 s 38976 0 39032 400 6 la_data_out[6]
port 176 nsew signal output
rlabel metal2 s 39648 0 39704 400 6 la_data_out[7]
port 177 nsew signal output
rlabel metal2 s 40320 0 40376 400 6 la_data_out[8]
port 178 nsew signal output
rlabel metal2 s 40992 0 41048 400 6 la_data_out[9]
port 179 nsew signal output
rlabel metal2 s 35168 0 35224 400 6 la_oenb[0]
port 180 nsew signal input
rlabel metal2 s 41888 0 41944 400 6 la_oenb[10]
port 181 nsew signal input
rlabel metal2 s 42560 0 42616 400 6 la_oenb[11]
port 182 nsew signal input
rlabel metal2 s 43232 0 43288 400 6 la_oenb[12]
port 183 nsew signal input
rlabel metal2 s 43904 0 43960 400 6 la_oenb[13]
port 184 nsew signal input
rlabel metal2 s 44576 0 44632 400 6 la_oenb[14]
port 185 nsew signal input
rlabel metal2 s 45248 0 45304 400 6 la_oenb[15]
port 186 nsew signal input
rlabel metal2 s 45920 0 45976 400 6 la_oenb[16]
port 187 nsew signal input
rlabel metal2 s 46592 0 46648 400 6 la_oenb[17]
port 188 nsew signal input
rlabel metal2 s 47264 0 47320 400 6 la_oenb[18]
port 189 nsew signal input
rlabel metal2 s 47936 0 47992 400 6 la_oenb[19]
port 190 nsew signal input
rlabel metal2 s 35840 0 35896 400 6 la_oenb[1]
port 191 nsew signal input
rlabel metal2 s 48608 0 48664 400 6 la_oenb[20]
port 192 nsew signal input
rlabel metal2 s 49280 0 49336 400 6 la_oenb[21]
port 193 nsew signal input
rlabel metal2 s 49952 0 50008 400 6 la_oenb[22]
port 194 nsew signal input
rlabel metal2 s 50624 0 50680 400 6 la_oenb[23]
port 195 nsew signal input
rlabel metal2 s 51296 0 51352 400 6 la_oenb[24]
port 196 nsew signal input
rlabel metal2 s 51968 0 52024 400 6 la_oenb[25]
port 197 nsew signal input
rlabel metal2 s 52640 0 52696 400 6 la_oenb[26]
port 198 nsew signal input
rlabel metal2 s 53312 0 53368 400 6 la_oenb[27]
port 199 nsew signal input
rlabel metal2 s 53984 0 54040 400 6 la_oenb[28]
port 200 nsew signal input
rlabel metal2 s 54656 0 54712 400 6 la_oenb[29]
port 201 nsew signal input
rlabel metal2 s 36512 0 36568 400 6 la_oenb[2]
port 202 nsew signal input
rlabel metal2 s 55328 0 55384 400 6 la_oenb[30]
port 203 nsew signal input
rlabel metal2 s 56000 0 56056 400 6 la_oenb[31]
port 204 nsew signal input
rlabel metal2 s 56672 0 56728 400 6 la_oenb[32]
port 205 nsew signal input
rlabel metal2 s 57344 0 57400 400 6 la_oenb[33]
port 206 nsew signal input
rlabel metal2 s 58016 0 58072 400 6 la_oenb[34]
port 207 nsew signal input
rlabel metal2 s 58688 0 58744 400 6 la_oenb[35]
port 208 nsew signal input
rlabel metal2 s 59360 0 59416 400 6 la_oenb[36]
port 209 nsew signal input
rlabel metal2 s 60032 0 60088 400 6 la_oenb[37]
port 210 nsew signal input
rlabel metal2 s 60704 0 60760 400 6 la_oenb[38]
port 211 nsew signal input
rlabel metal2 s 61376 0 61432 400 6 la_oenb[39]
port 212 nsew signal input
rlabel metal2 s 37184 0 37240 400 6 la_oenb[3]
port 213 nsew signal input
rlabel metal2 s 62048 0 62104 400 6 la_oenb[40]
port 214 nsew signal input
rlabel metal2 s 62720 0 62776 400 6 la_oenb[41]
port 215 nsew signal input
rlabel metal2 s 63392 0 63448 400 6 la_oenb[42]
port 216 nsew signal input
rlabel metal2 s 64064 0 64120 400 6 la_oenb[43]
port 217 nsew signal input
rlabel metal2 s 64736 0 64792 400 6 la_oenb[44]
port 218 nsew signal input
rlabel metal2 s 65408 0 65464 400 6 la_oenb[45]
port 219 nsew signal input
rlabel metal2 s 66080 0 66136 400 6 la_oenb[46]
port 220 nsew signal input
rlabel metal2 s 66752 0 66808 400 6 la_oenb[47]
port 221 nsew signal input
rlabel metal2 s 67424 0 67480 400 6 la_oenb[48]
port 222 nsew signal input
rlabel metal2 s 68096 0 68152 400 6 la_oenb[49]
port 223 nsew signal input
rlabel metal2 s 37856 0 37912 400 6 la_oenb[4]
port 224 nsew signal input
rlabel metal2 s 68768 0 68824 400 6 la_oenb[50]
port 225 nsew signal input
rlabel metal2 s 69440 0 69496 400 6 la_oenb[51]
port 226 nsew signal input
rlabel metal2 s 70112 0 70168 400 6 la_oenb[52]
port 227 nsew signal input
rlabel metal2 s 70784 0 70840 400 6 la_oenb[53]
port 228 nsew signal input
rlabel metal2 s 71456 0 71512 400 6 la_oenb[54]
port 229 nsew signal input
rlabel metal2 s 72128 0 72184 400 6 la_oenb[55]
port 230 nsew signal input
rlabel metal2 s 72800 0 72856 400 6 la_oenb[56]
port 231 nsew signal input
rlabel metal2 s 73472 0 73528 400 6 la_oenb[57]
port 232 nsew signal input
rlabel metal2 s 74144 0 74200 400 6 la_oenb[58]
port 233 nsew signal input
rlabel metal2 s 74816 0 74872 400 6 la_oenb[59]
port 234 nsew signal input
rlabel metal2 s 38528 0 38584 400 6 la_oenb[5]
port 235 nsew signal input
rlabel metal2 s 75488 0 75544 400 6 la_oenb[60]
port 236 nsew signal input
rlabel metal2 s 76160 0 76216 400 6 la_oenb[61]
port 237 nsew signal input
rlabel metal2 s 76832 0 76888 400 6 la_oenb[62]
port 238 nsew signal input
rlabel metal2 s 77504 0 77560 400 6 la_oenb[63]
port 239 nsew signal input
rlabel metal2 s 39200 0 39256 400 6 la_oenb[6]
port 240 nsew signal input
rlabel metal2 s 39872 0 39928 400 6 la_oenb[7]
port 241 nsew signal input
rlabel metal2 s 40544 0 40600 400 6 la_oenb[8]
port 242 nsew signal input
rlabel metal2 s 41216 0 41272 400 6 la_oenb[9]
port 243 nsew signal input
rlabel metal4 s 2224 1538 2384 89406 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 89406 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 89406 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 89406 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 89406 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 89406 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 89406 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 89406 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 89406 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 89406 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 89406 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 89406 6 vss
port 245 nsew ground bidirectional
rlabel metal2 s 10976 0 11032 400 6 wb_clk_i
port 246 nsew signal input
rlabel metal2 s 11200 0 11256 400 6 wb_rst_i
port 247 nsew signal input
rlabel metal2 s 11424 0 11480 400 6 wbs_ack_o
port 248 nsew signal output
rlabel metal2 s 12320 0 12376 400 6 wbs_adr_i[0]
port 249 nsew signal input
rlabel metal2 s 19936 0 19992 400 6 wbs_adr_i[10]
port 250 nsew signal input
rlabel metal2 s 20608 0 20664 400 6 wbs_adr_i[11]
port 251 nsew signal input
rlabel metal2 s 21280 0 21336 400 6 wbs_adr_i[12]
port 252 nsew signal input
rlabel metal2 s 21952 0 22008 400 6 wbs_adr_i[13]
port 253 nsew signal input
rlabel metal2 s 22624 0 22680 400 6 wbs_adr_i[14]
port 254 nsew signal input
rlabel metal2 s 23296 0 23352 400 6 wbs_adr_i[15]
port 255 nsew signal input
rlabel metal2 s 23968 0 24024 400 6 wbs_adr_i[16]
port 256 nsew signal input
rlabel metal2 s 24640 0 24696 400 6 wbs_adr_i[17]
port 257 nsew signal input
rlabel metal2 s 25312 0 25368 400 6 wbs_adr_i[18]
port 258 nsew signal input
rlabel metal2 s 25984 0 26040 400 6 wbs_adr_i[19]
port 259 nsew signal input
rlabel metal2 s 13216 0 13272 400 6 wbs_adr_i[1]
port 260 nsew signal input
rlabel metal2 s 26656 0 26712 400 6 wbs_adr_i[20]
port 261 nsew signal input
rlabel metal2 s 27328 0 27384 400 6 wbs_adr_i[21]
port 262 nsew signal input
rlabel metal2 s 28000 0 28056 400 6 wbs_adr_i[22]
port 263 nsew signal input
rlabel metal2 s 28672 0 28728 400 6 wbs_adr_i[23]
port 264 nsew signal input
rlabel metal2 s 29344 0 29400 400 6 wbs_adr_i[24]
port 265 nsew signal input
rlabel metal2 s 30016 0 30072 400 6 wbs_adr_i[25]
port 266 nsew signal input
rlabel metal2 s 30688 0 30744 400 6 wbs_adr_i[26]
port 267 nsew signal input
rlabel metal2 s 31360 0 31416 400 6 wbs_adr_i[27]
port 268 nsew signal input
rlabel metal2 s 32032 0 32088 400 6 wbs_adr_i[28]
port 269 nsew signal input
rlabel metal2 s 32704 0 32760 400 6 wbs_adr_i[29]
port 270 nsew signal input
rlabel metal2 s 14112 0 14168 400 6 wbs_adr_i[2]
port 271 nsew signal input
rlabel metal2 s 33376 0 33432 400 6 wbs_adr_i[30]
port 272 nsew signal input
rlabel metal2 s 34048 0 34104 400 6 wbs_adr_i[31]
port 273 nsew signal input
rlabel metal2 s 15008 0 15064 400 6 wbs_adr_i[3]
port 274 nsew signal input
rlabel metal2 s 15904 0 15960 400 6 wbs_adr_i[4]
port 275 nsew signal input
rlabel metal2 s 16576 0 16632 400 6 wbs_adr_i[5]
port 276 nsew signal input
rlabel metal2 s 17248 0 17304 400 6 wbs_adr_i[6]
port 277 nsew signal input
rlabel metal2 s 17920 0 17976 400 6 wbs_adr_i[7]
port 278 nsew signal input
rlabel metal2 s 18592 0 18648 400 6 wbs_adr_i[8]
port 279 nsew signal input
rlabel metal2 s 19264 0 19320 400 6 wbs_adr_i[9]
port 280 nsew signal input
rlabel metal2 s 11648 0 11704 400 6 wbs_cyc_i
port 281 nsew signal input
rlabel metal2 s 12544 0 12600 400 6 wbs_dat_i[0]
port 282 nsew signal input
rlabel metal2 s 20160 0 20216 400 6 wbs_dat_i[10]
port 283 nsew signal input
rlabel metal2 s 20832 0 20888 400 6 wbs_dat_i[11]
port 284 nsew signal input
rlabel metal2 s 21504 0 21560 400 6 wbs_dat_i[12]
port 285 nsew signal input
rlabel metal2 s 22176 0 22232 400 6 wbs_dat_i[13]
port 286 nsew signal input
rlabel metal2 s 22848 0 22904 400 6 wbs_dat_i[14]
port 287 nsew signal input
rlabel metal2 s 23520 0 23576 400 6 wbs_dat_i[15]
port 288 nsew signal input
rlabel metal2 s 24192 0 24248 400 6 wbs_dat_i[16]
port 289 nsew signal input
rlabel metal2 s 24864 0 24920 400 6 wbs_dat_i[17]
port 290 nsew signal input
rlabel metal2 s 25536 0 25592 400 6 wbs_dat_i[18]
port 291 nsew signal input
rlabel metal2 s 26208 0 26264 400 6 wbs_dat_i[19]
port 292 nsew signal input
rlabel metal2 s 13440 0 13496 400 6 wbs_dat_i[1]
port 293 nsew signal input
rlabel metal2 s 26880 0 26936 400 6 wbs_dat_i[20]
port 294 nsew signal input
rlabel metal2 s 27552 0 27608 400 6 wbs_dat_i[21]
port 295 nsew signal input
rlabel metal2 s 28224 0 28280 400 6 wbs_dat_i[22]
port 296 nsew signal input
rlabel metal2 s 28896 0 28952 400 6 wbs_dat_i[23]
port 297 nsew signal input
rlabel metal2 s 29568 0 29624 400 6 wbs_dat_i[24]
port 298 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 wbs_dat_i[25]
port 299 nsew signal input
rlabel metal2 s 30912 0 30968 400 6 wbs_dat_i[26]
port 300 nsew signal input
rlabel metal2 s 31584 0 31640 400 6 wbs_dat_i[27]
port 301 nsew signal input
rlabel metal2 s 32256 0 32312 400 6 wbs_dat_i[28]
port 302 nsew signal input
rlabel metal2 s 32928 0 32984 400 6 wbs_dat_i[29]
port 303 nsew signal input
rlabel metal2 s 14336 0 14392 400 6 wbs_dat_i[2]
port 304 nsew signal input
rlabel metal2 s 33600 0 33656 400 6 wbs_dat_i[30]
port 305 nsew signal input
rlabel metal2 s 34272 0 34328 400 6 wbs_dat_i[31]
port 306 nsew signal input
rlabel metal2 s 15232 0 15288 400 6 wbs_dat_i[3]
port 307 nsew signal input
rlabel metal2 s 16128 0 16184 400 6 wbs_dat_i[4]
port 308 nsew signal input
rlabel metal2 s 16800 0 16856 400 6 wbs_dat_i[5]
port 309 nsew signal input
rlabel metal2 s 17472 0 17528 400 6 wbs_dat_i[6]
port 310 nsew signal input
rlabel metal2 s 18144 0 18200 400 6 wbs_dat_i[7]
port 311 nsew signal input
rlabel metal2 s 18816 0 18872 400 6 wbs_dat_i[8]
port 312 nsew signal input
rlabel metal2 s 19488 0 19544 400 6 wbs_dat_i[9]
port 313 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 wbs_dat_o[0]
port 314 nsew signal output
rlabel metal2 s 20384 0 20440 400 6 wbs_dat_o[10]
port 315 nsew signal output
rlabel metal2 s 21056 0 21112 400 6 wbs_dat_o[11]
port 316 nsew signal output
rlabel metal2 s 21728 0 21784 400 6 wbs_dat_o[12]
port 317 nsew signal output
rlabel metal2 s 22400 0 22456 400 6 wbs_dat_o[13]
port 318 nsew signal output
rlabel metal2 s 23072 0 23128 400 6 wbs_dat_o[14]
port 319 nsew signal output
rlabel metal2 s 23744 0 23800 400 6 wbs_dat_o[15]
port 320 nsew signal output
rlabel metal2 s 24416 0 24472 400 6 wbs_dat_o[16]
port 321 nsew signal output
rlabel metal2 s 25088 0 25144 400 6 wbs_dat_o[17]
port 322 nsew signal output
rlabel metal2 s 25760 0 25816 400 6 wbs_dat_o[18]
port 323 nsew signal output
rlabel metal2 s 26432 0 26488 400 6 wbs_dat_o[19]
port 324 nsew signal output
rlabel metal2 s 13664 0 13720 400 6 wbs_dat_o[1]
port 325 nsew signal output
rlabel metal2 s 27104 0 27160 400 6 wbs_dat_o[20]
port 326 nsew signal output
rlabel metal2 s 27776 0 27832 400 6 wbs_dat_o[21]
port 327 nsew signal output
rlabel metal2 s 28448 0 28504 400 6 wbs_dat_o[22]
port 328 nsew signal output
rlabel metal2 s 29120 0 29176 400 6 wbs_dat_o[23]
port 329 nsew signal output
rlabel metal2 s 29792 0 29848 400 6 wbs_dat_o[24]
port 330 nsew signal output
rlabel metal2 s 30464 0 30520 400 6 wbs_dat_o[25]
port 331 nsew signal output
rlabel metal2 s 31136 0 31192 400 6 wbs_dat_o[26]
port 332 nsew signal output
rlabel metal2 s 31808 0 31864 400 6 wbs_dat_o[27]
port 333 nsew signal output
rlabel metal2 s 32480 0 32536 400 6 wbs_dat_o[28]
port 334 nsew signal output
rlabel metal2 s 33152 0 33208 400 6 wbs_dat_o[29]
port 335 nsew signal output
rlabel metal2 s 14560 0 14616 400 6 wbs_dat_o[2]
port 336 nsew signal output
rlabel metal2 s 33824 0 33880 400 6 wbs_dat_o[30]
port 337 nsew signal output
rlabel metal2 s 34496 0 34552 400 6 wbs_dat_o[31]
port 338 nsew signal output
rlabel metal2 s 15456 0 15512 400 6 wbs_dat_o[3]
port 339 nsew signal output
rlabel metal2 s 16352 0 16408 400 6 wbs_dat_o[4]
port 340 nsew signal output
rlabel metal2 s 17024 0 17080 400 6 wbs_dat_o[5]
port 341 nsew signal output
rlabel metal2 s 17696 0 17752 400 6 wbs_dat_o[6]
port 342 nsew signal output
rlabel metal2 s 18368 0 18424 400 6 wbs_dat_o[7]
port 343 nsew signal output
rlabel metal2 s 19040 0 19096 400 6 wbs_dat_o[8]
port 344 nsew signal output
rlabel metal2 s 19712 0 19768 400 6 wbs_dat_o[9]
port 345 nsew signal output
rlabel metal2 s 12992 0 13048 400 6 wbs_sel_i[0]
port 346 nsew signal input
rlabel metal2 s 13888 0 13944 400 6 wbs_sel_i[1]
port 347 nsew signal input
rlabel metal2 s 14784 0 14840 400 6 wbs_sel_i[2]
port 348 nsew signal input
rlabel metal2 s 15680 0 15736 400 6 wbs_sel_i[3]
port 349 nsew signal input
rlabel metal2 s 11872 0 11928 400 6 wbs_stb_i
port 350 nsew signal input
rlabel metal2 s 12096 0 12152 400 6 wbs_we_i
port 351 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 89371 91163
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 23964264
string GDS_FILE /home/kris/repos/diy-ic/lincoln-gfmpw-1d/openlane/user_proj_example/runs/23_12_07_21_03/results/signoff/user_proj_example.magic.gds
string GDS_START 520002
<< end >>

