VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ram_6x64
  CLASS BLOCK ;
  FOREIGN ram_6x64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 777.420 BY 795.340 ;
  PIN address_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 773.420 440.160 777.420 440.720 ;
    END
  END address_i[0]
  PIN address_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 773.420 231.840 777.420 232.400 ;
    END
  END address_i[1]
  PIN address_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 773.420 322.560 777.420 323.120 ;
    END
  END address_i[2]
  PIN address_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 0.000 363.440 4.000 ;
    END
  END address_i[3]
  PIN address_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 0.000 366.800 4.000 ;
    END
  END address_i[4]
  PIN address_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 0.000 370.160 4.000 ;
    END
  END address_i[5]
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 766.080 4.000 766.640 ;
    END
  END clk_i
  PIN data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 0.000 339.920 4.000 ;
    END
  END data_i[0]
  PIN data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 773.420 426.720 777.420 427.280 ;
    END
  END data_i[10]
  PIN data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 773.420 433.440 777.420 434.000 ;
    END
  END data_i[11]
  PIN data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 773.420 443.520 777.420 444.080 ;
    END
  END data_i[12]
  PIN data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 773.420 450.240 777.420 450.800 ;
    END
  END data_i[13]
  PIN data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 791.340 487.760 795.340 ;
    END
  END data_i[14]
  PIN data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 791.340 477.680 795.340 ;
    END
  END data_i[15]
  PIN data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 791.340 481.040 795.340 ;
    END
  END data_i[16]
  PIN data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 791.340 484.400 795.340 ;
    END
  END data_i[17]
  PIN data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 791.340 491.120 795.340 ;
    END
  END data_i[18]
  PIN data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 791.340 494.480 795.340 ;
    END
  END data_i[19]
  PIN data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 0.000 329.840 4.000 ;
    END
  END data_i[1]
  PIN data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 456.960 4.000 457.520 ;
    END
  END data_i[20]
  PIN data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 460.320 4.000 460.880 ;
    END
  END data_i[21]
  PIN data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 483.840 4.000 484.400 ;
    END
  END data_i[22]
  PIN data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 463.680 4.000 464.240 ;
    END
  END data_i[23]
  PIN data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 470.400 4.000 470.960 ;
    END
  END data_i[24]
  PIN data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 473.760 4.000 474.320 ;
    END
  END data_i[25]
  PIN data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 490.560 4.000 491.120 ;
    END
  END data_i[26]
  PIN data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 480.480 4.000 481.040 ;
    END
  END data_i[27]
  PIN data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 467.040 4.000 467.600 ;
    END
  END data_i[28]
  PIN data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 487.200 4.000 487.760 ;
    END
  END data_i[29]
  PIN data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 0.000 313.040 4.000 ;
    END
  END data_i[2]
  PIN data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 0.000 286.160 4.000 ;
    END
  END data_i[30]
  PIN data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 0.000 289.520 4.000 ;
    END
  END data_i[31]
  PIN data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 0.000 333.200 4.000 ;
    END
  END data_i[3]
  PIN data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 0.000 323.120 4.000 ;
    END
  END data_i[4]
  PIN data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 0.000 306.320 4.000 ;
    END
  END data_i[5]
  PIN data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 0.000 309.680 4.000 ;
    END
  END data_i[6]
  PIN data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 0.000 299.600 4.000 ;
    END
  END data_i[7]
  PIN data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 0.000 292.880 4.000 ;
    END
  END data_i[8]
  PIN data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 0.000 302.960 4.000 ;
    END
  END data_i[9]
  PIN data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 0.000 497.840 4.000 ;
    END
  END data_o[0]
  PIN data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 773.420 460.320 777.420 460.880 ;
    END
  END data_o[10]
  PIN data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 791.340 507.920 795.340 ;
    END
  END data_o[11]
  PIN data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 773.420 456.960 777.420 457.520 ;
    END
  END data_o[12]
  PIN data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 791.340 504.560 795.340 ;
    END
  END data_o[13]
  PIN data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 773.420 477.120 777.420 477.680 ;
    END
  END data_o[14]
  PIN data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 773.420 473.760 777.420 474.320 ;
    END
  END data_o[15]
  PIN data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 791.340 521.360 795.340 ;
    END
  END data_o[16]
  PIN data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 791.340 501.200 795.340 ;
    END
  END data_o[17]
  PIN data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 791.340 511.280 795.340 ;
    END
  END data_o[18]
  PIN data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 791.340 497.840 795.340 ;
    END
  END data_o[19]
  PIN data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 0.000 494.480 4.000 ;
    END
  END data_o[1]
  PIN data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 571.200 4.000 571.760 ;
    END
  END data_o[20]
  PIN data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 574.560 4.000 575.120 ;
    END
  END data_o[21]
  PIN data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 554.400 4.000 554.960 ;
    END
  END data_o[22]
  PIN data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 567.840 4.000 568.400 ;
    END
  END data_o[23]
  PIN data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 534.240 4.000 534.800 ;
    END
  END data_o[24]
  PIN data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 544.320 4.000 544.880 ;
    END
  END data_o[25]
  PIN data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 520.800 4.000 521.360 ;
    END
  END data_o[26]
  PIN data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 504.000 4.000 504.560 ;
    END
  END data_o[27]
  PIN data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 493.920 4.000 494.480 ;
    END
  END data_o[28]
  PIN data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 477.120 4.000 477.680 ;
    END
  END data_o[29]
  PIN data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 0.000 501.200 4.000 ;
    END
  END data_o[2]
  PIN data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 265.440 4.000 266.000 ;
    END
  END data_o[30]
  PIN data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.080 4.000 262.640 ;
    END
  END data_o[31]
  PIN data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 0.000 504.560 4.000 ;
    END
  END data_o[3]
  PIN data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 0.000 689.360 4.000 ;
    END
  END data_o[4]
  PIN data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 675.360 0.000 675.920 4.000 ;
    END
  END data_o[5]
  PIN data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 0.000 682.640 4.000 ;
    END
  END data_o[6]
  PIN data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 0.000 679.280 4.000 ;
    END
  END data_o[7]
  PIN data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 0.000 672.560 4.000 ;
    END
  END data_o[8]
  PIN data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 0.000 686.000 4.000 ;
    END
  END data_o[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 776.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 776.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 776.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 776.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 776.460 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 776.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 776.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 776.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 776.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 776.460 ;
    END
  END vss
  PIN we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 770.560 777.690 ;
      LAYER Metal2 ;
        RECT 0.140 791.040 476.820 791.340 ;
        RECT 477.980 791.040 480.180 791.340 ;
        RECT 481.340 791.040 483.540 791.340 ;
        RECT 484.700 791.040 486.900 791.340 ;
        RECT 488.060 791.040 490.260 791.340 ;
        RECT 491.420 791.040 493.620 791.340 ;
        RECT 494.780 791.040 496.980 791.340 ;
        RECT 498.140 791.040 500.340 791.340 ;
        RECT 501.500 791.040 503.700 791.340 ;
        RECT 504.860 791.040 507.060 791.340 ;
        RECT 508.220 791.040 510.420 791.340 ;
        RECT 511.580 791.040 520.500 791.340 ;
        RECT 521.660 791.040 768.740 791.340 ;
        RECT 0.140 4.300 768.740 791.040 ;
        RECT 0.140 3.500 285.300 4.300 ;
        RECT 286.460 3.500 288.660 4.300 ;
        RECT 289.820 3.500 292.020 4.300 ;
        RECT 293.180 3.500 298.740 4.300 ;
        RECT 299.900 3.500 302.100 4.300 ;
        RECT 303.260 3.500 305.460 4.300 ;
        RECT 306.620 3.500 308.820 4.300 ;
        RECT 309.980 3.500 312.180 4.300 ;
        RECT 313.340 3.500 322.260 4.300 ;
        RECT 323.420 3.500 328.980 4.300 ;
        RECT 330.140 3.500 332.340 4.300 ;
        RECT 333.500 3.500 339.060 4.300 ;
        RECT 340.220 3.500 362.580 4.300 ;
        RECT 363.740 3.500 365.940 4.300 ;
        RECT 367.100 3.500 369.300 4.300 ;
        RECT 370.460 3.500 493.620 4.300 ;
        RECT 494.780 3.500 496.980 4.300 ;
        RECT 498.140 3.500 500.340 4.300 ;
        RECT 501.500 3.500 503.700 4.300 ;
        RECT 504.860 3.500 671.700 4.300 ;
        RECT 672.860 3.500 675.060 4.300 ;
        RECT 676.220 3.500 678.420 4.300 ;
        RECT 679.580 3.500 681.780 4.300 ;
        RECT 682.940 3.500 685.140 4.300 ;
        RECT 686.300 3.500 688.500 4.300 ;
        RECT 689.660 3.500 768.740 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 766.940 773.420 776.300 ;
        RECT 4.300 765.780 773.420 766.940 ;
        RECT 0.090 575.420 773.420 765.780 ;
        RECT 4.300 574.260 773.420 575.420 ;
        RECT 0.090 572.060 773.420 574.260 ;
        RECT 4.300 570.900 773.420 572.060 ;
        RECT 0.090 568.700 773.420 570.900 ;
        RECT 4.300 567.540 773.420 568.700 ;
        RECT 0.090 555.260 773.420 567.540 ;
        RECT 4.300 554.100 773.420 555.260 ;
        RECT 0.090 545.180 773.420 554.100 ;
        RECT 4.300 544.020 773.420 545.180 ;
        RECT 0.090 535.100 773.420 544.020 ;
        RECT 4.300 533.940 773.420 535.100 ;
        RECT 0.090 521.660 773.420 533.940 ;
        RECT 4.300 520.500 773.420 521.660 ;
        RECT 0.090 504.860 773.420 520.500 ;
        RECT 4.300 503.700 773.420 504.860 ;
        RECT 0.090 494.780 773.420 503.700 ;
        RECT 4.300 493.620 773.420 494.780 ;
        RECT 0.090 491.420 773.420 493.620 ;
        RECT 4.300 490.260 773.420 491.420 ;
        RECT 0.090 488.060 773.420 490.260 ;
        RECT 4.300 486.900 773.420 488.060 ;
        RECT 0.090 484.700 773.420 486.900 ;
        RECT 4.300 483.540 773.420 484.700 ;
        RECT 0.090 481.340 773.420 483.540 ;
        RECT 4.300 480.180 773.420 481.340 ;
        RECT 0.090 477.980 773.420 480.180 ;
        RECT 4.300 476.820 773.120 477.980 ;
        RECT 0.090 474.620 773.420 476.820 ;
        RECT 4.300 473.460 773.120 474.620 ;
        RECT 0.090 471.260 773.420 473.460 ;
        RECT 4.300 470.100 773.420 471.260 ;
        RECT 0.090 467.900 773.420 470.100 ;
        RECT 4.300 466.740 773.420 467.900 ;
        RECT 0.090 464.540 773.420 466.740 ;
        RECT 4.300 463.380 773.420 464.540 ;
        RECT 0.090 461.180 773.420 463.380 ;
        RECT 4.300 460.020 773.120 461.180 ;
        RECT 0.090 457.820 773.420 460.020 ;
        RECT 4.300 456.660 773.120 457.820 ;
        RECT 0.090 451.100 773.420 456.660 ;
        RECT 0.090 449.940 773.120 451.100 ;
        RECT 0.090 444.380 773.420 449.940 ;
        RECT 0.090 443.220 773.120 444.380 ;
        RECT 0.090 441.020 773.420 443.220 ;
        RECT 0.090 439.860 773.120 441.020 ;
        RECT 0.090 434.300 773.420 439.860 ;
        RECT 0.090 433.140 773.120 434.300 ;
        RECT 0.090 427.580 773.420 433.140 ;
        RECT 0.090 426.420 773.120 427.580 ;
        RECT 0.090 323.420 773.420 426.420 ;
        RECT 0.090 322.260 773.120 323.420 ;
        RECT 0.090 266.300 773.420 322.260 ;
        RECT 4.300 265.140 773.420 266.300 ;
        RECT 0.090 262.940 773.420 265.140 ;
        RECT 4.300 261.780 773.420 262.940 ;
        RECT 0.090 232.700 773.420 261.780 ;
        RECT 0.090 231.540 773.120 232.700 ;
        RECT 0.090 121.820 773.420 231.540 ;
        RECT 4.300 120.660 773.420 121.820 ;
        RECT 0.090 6.300 773.420 120.660 ;
      LAYER Metal4 ;
        RECT 56.700 16.890 98.740 773.830 ;
        RECT 100.940 16.890 175.540 773.830 ;
        RECT 177.740 16.890 252.340 773.830 ;
        RECT 254.540 16.890 329.140 773.830 ;
        RECT 331.340 16.890 405.940 773.830 ;
        RECT 408.140 16.890 482.740 773.830 ;
        RECT 484.940 16.890 559.540 773.830 ;
        RECT 561.740 16.890 636.340 773.830 ;
        RECT 638.540 16.890 713.140 773.830 ;
        RECT 715.340 16.890 722.260 773.830 ;
  END
END ram_6x64
END LIBRARY

