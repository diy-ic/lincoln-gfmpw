magic
tech gf180mcuD
magscale 1 5
timestamp 1701783335
<< obsm1 >>
rect 672 1471 9455 8385
<< metal2 >>
rect 0 9600 56 10000
rect 336 9600 392 10000
rect 672 9600 728 10000
rect 1008 9600 1064 10000
rect 1344 9600 1400 10000
rect 1680 9600 1736 10000
rect 2016 9600 2072 10000
rect 2352 9600 2408 10000
rect 2688 9600 2744 10000
rect 3024 9600 3080 10000
rect 3360 9600 3416 10000
rect 3696 9600 3752 10000
rect 4032 9600 4088 10000
rect 4368 9600 4424 10000
rect 4704 9600 4760 10000
rect 5040 9600 5096 10000
rect 5376 9600 5432 10000
rect 5712 9600 5768 10000
rect 6048 9600 6104 10000
rect 6384 9600 6440 10000
rect 6720 9600 6776 10000
rect 7056 9600 7112 10000
rect 7392 9600 7448 10000
rect 7728 9600 7784 10000
rect 8064 9600 8120 10000
rect 8400 9600 8456 10000
rect 8736 9600 8792 10000
rect 9072 9600 9128 10000
rect 9408 9600 9464 10000
rect 9744 9600 9800 10000
rect 0 0 56 400
rect 336 0 392 400
rect 672 0 728 400
rect 1008 0 1064 400
rect 1344 0 1400 400
rect 1680 0 1736 400
rect 2016 0 2072 400
rect 2352 0 2408 400
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 4032 0 4088 400
rect 4368 0 4424 400
rect 4704 0 4760 400
rect 5040 0 5096 400
rect 5376 0 5432 400
rect 5712 0 5768 400
rect 6048 0 6104 400
rect 6384 0 6440 400
rect 6720 0 6776 400
rect 7056 0 7112 400
rect 7392 0 7448 400
rect 7728 0 7784 400
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 9744 0 9800 400
<< obsm2 >>
rect 86 9570 306 9600
rect 422 9570 642 9600
rect 758 9570 978 9600
rect 1094 9570 1314 9600
rect 1430 9570 1650 9600
rect 1766 9570 1986 9600
rect 2102 9570 2322 9600
rect 2438 9570 2658 9600
rect 2774 9570 2994 9600
rect 3110 9570 3330 9600
rect 3446 9570 3666 9600
rect 3782 9570 4002 9600
rect 4118 9570 4338 9600
rect 4454 9570 4674 9600
rect 4790 9570 5010 9600
rect 5126 9570 5346 9600
rect 5462 9570 5682 9600
rect 5798 9570 6018 9600
rect 6134 9570 6354 9600
rect 6470 9570 6690 9600
rect 6806 9570 7026 9600
rect 7142 9570 7362 9600
rect 7478 9570 7698 9600
rect 7814 9570 8034 9600
rect 8150 9570 8370 9600
rect 8486 9570 8706 9600
rect 8822 9570 9042 9600
rect 9158 9570 9378 9600
rect 9494 9570 9714 9600
rect 14 430 9786 9570
rect 86 400 306 430
rect 422 400 642 430
rect 758 400 978 430
rect 1094 400 1314 430
rect 1430 400 1650 430
rect 1766 400 1986 430
rect 2102 400 2322 430
rect 2438 400 2658 430
rect 2774 400 2994 430
rect 3110 400 3330 430
rect 3446 400 3666 430
rect 3782 400 4002 430
rect 4118 400 4338 430
rect 4454 400 4674 430
rect 4790 400 5010 430
rect 5126 400 5346 430
rect 5462 400 5682 430
rect 5798 400 6018 430
rect 6134 400 6354 430
rect 6470 400 6690 430
rect 6806 400 7026 430
rect 7142 400 7362 430
rect 7478 400 7698 430
rect 7814 400 8034 430
rect 8150 400 8370 430
rect 8486 400 8706 430
rect 8822 400 9042 430
rect 9158 400 9378 430
rect 9494 400 9714 430
<< metal3 >>
rect 0 9744 400 9800
rect 9600 9744 10000 9800
rect 0 9408 400 9464
rect 9600 9408 10000 9464
rect 0 9072 400 9128
rect 9600 9072 10000 9128
rect 0 8736 400 8792
rect 9600 8736 10000 8792
rect 9600 8400 10000 8456
rect 9600 8064 10000 8120
rect 0 7728 400 7784
rect 9600 7728 10000 7784
rect 0 7392 400 7448
rect 9600 7392 10000 7448
rect 0 7056 400 7112
rect 9600 7056 10000 7112
rect 0 6720 400 6776
rect 9600 6720 10000 6776
rect 9600 6384 10000 6440
rect 0 6048 400 6104
rect 9600 6048 10000 6104
rect 0 5712 400 5768
rect 9600 5712 10000 5768
rect 0 5376 400 5432
rect 9600 5376 10000 5432
rect 0 5040 400 5096
rect 9600 5040 10000 5096
rect 9600 4704 10000 4760
rect 9600 4368 10000 4424
rect 0 4032 400 4088
rect 9600 4032 10000 4088
rect 0 3696 400 3752
rect 9600 3696 10000 3752
rect 9600 3360 10000 3416
rect 9600 3024 10000 3080
rect 0 2688 400 2744
rect 9600 2688 10000 2744
rect 0 2352 400 2408
rect 9600 2352 10000 2408
rect 0 2016 400 2072
rect 9600 2016 10000 2072
rect 9600 1680 10000 1736
rect 9600 1344 10000 1400
rect 9600 1008 10000 1064
rect 9600 672 10000 728
rect 9600 336 10000 392
rect 9600 0 10000 56
<< obsm3 >>
rect 9 8150 9791 8246
rect 9 8034 9570 8150
rect 9 7814 9791 8034
rect 430 7698 9570 7814
rect 9 7478 9791 7698
rect 430 7362 9570 7478
rect 9 7142 9791 7362
rect 430 7026 9570 7142
rect 9 6806 9791 7026
rect 430 6690 9570 6806
rect 9 6470 9791 6690
rect 9 6354 9570 6470
rect 9 6134 9791 6354
rect 430 6018 9570 6134
rect 9 5798 9791 6018
rect 430 5682 9570 5798
rect 9 5462 9791 5682
rect 430 5346 9570 5462
rect 9 5126 9791 5346
rect 430 5010 9570 5126
rect 9 4790 9791 5010
rect 9 4674 9570 4790
rect 9 4454 9791 4674
rect 9 4338 9570 4454
rect 9 4118 9791 4338
rect 430 4002 9570 4118
rect 9 3782 9791 4002
rect 430 3666 9570 3782
rect 9 3446 9791 3666
rect 9 3330 9570 3446
rect 9 3110 9791 3330
rect 9 2994 9570 3110
rect 9 2774 9791 2994
rect 430 2658 9570 2774
rect 9 2438 9791 2658
rect 430 2322 9570 2438
rect 9 2102 9791 2322
rect 430 1986 9570 2102
rect 9 1766 9791 1986
rect 9 1650 9570 1766
rect 9 1554 9791 1650
<< metal4 >>
rect 1670 1538 1830 8262
rect 2748 1538 2908 8262
rect 3826 1538 3986 8262
rect 4904 1538 5064 8262
rect 5982 1538 6142 8262
rect 7060 1538 7220 8262
rect 8138 1538 8298 8262
rect 9216 1538 9376 8262
<< labels >>
rlabel metal2 s 1344 9600 1400 10000 6 reg_q_o
port 1 nsew signal output
rlabel metal4 s 1670 1538 1830 8262 6 vdd
port 2 nsew power bidirectional
rlabel metal4 s 3826 1538 3986 8262 6 vdd
port 2 nsew power bidirectional
rlabel metal4 s 5982 1538 6142 8262 6 vdd
port 2 nsew power bidirectional
rlabel metal4 s 8138 1538 8298 8262 6 vdd
port 2 nsew power bidirectional
rlabel metal4 s 2748 1538 2908 8262 6 vss
port 3 nsew ground bidirectional
rlabel metal4 s 4904 1538 5064 8262 6 vss
port 3 nsew ground bidirectional
rlabel metal4 s 7060 1538 7220 8262 6 vss
port 3 nsew ground bidirectional
rlabel metal4 s 9216 1538 9376 8262 6 vss
port 3 nsew ground bidirectional
rlabel metal3 s 0 6048 400 6104 6 wb_clk_i
port 4 nsew signal input
rlabel metal2 s 3696 9600 3752 10000 6 wb_rst_i
port 5 nsew signal input
rlabel metal2 s 2352 9600 2408 10000 6 wbs_ack_o
port 6 nsew signal output
rlabel metal2 s 9408 0 9464 400 6 wbs_adr_i[0]
port 7 nsew signal input
rlabel metal2 s 0 0 56 400 6 wbs_adr_i[10]
port 8 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 wbs_adr_i[11]
port 9 nsew signal input
rlabel metal2 s 336 0 392 400 6 wbs_adr_i[12]
port 10 nsew signal input
rlabel metal2 s 672 0 728 400 6 wbs_adr_i[13]
port 11 nsew signal input
rlabel metal2 s 1680 0 1736 400 6 wbs_adr_i[14]
port 12 nsew signal input
rlabel metal2 s 1344 0 1400 400 6 wbs_adr_i[15]
port 13 nsew signal input
rlabel metal2 s 2352 0 2408 400 6 wbs_adr_i[16]
port 14 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 wbs_adr_i[17]
port 15 nsew signal input
rlabel metal2 s 2688 0 2744 400 6 wbs_adr_i[18]
port 16 nsew signal input
rlabel metal2 s 2016 0 2072 400 6 wbs_adr_i[19]
port 17 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 wbs_adr_i[1]
port 18 nsew signal input
rlabel metal2 s 4032 0 4088 400 6 wbs_adr_i[20]
port 19 nsew signal input
rlabel metal2 s 3696 0 3752 400 6 wbs_adr_i[21]
port 20 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 wbs_adr_i[22]
port 21 nsew signal input
rlabel metal3 s 9600 4368 10000 4424 6 wbs_adr_i[23]
port 22 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 wbs_adr_i[24]
port 23 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 wbs_adr_i[25]
port 24 nsew signal input
rlabel metal2 s 6384 0 6440 400 6 wbs_adr_i[26]
port 25 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 wbs_adr_i[27]
port 26 nsew signal input
rlabel metal3 s 9600 3696 10000 3752 6 wbs_adr_i[28]
port 27 nsew signal input
rlabel metal3 s 9600 4032 10000 4088 6 wbs_adr_i[29]
port 28 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 wbs_adr_i[2]
port 29 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 wbs_adr_i[30]
port 30 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 wbs_adr_i[31]
port 31 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 wbs_adr_i[3]
port 32 nsew signal input
rlabel metal2 s 5376 0 5432 400 6 wbs_adr_i[4]
port 33 nsew signal input
rlabel metal2 s 5712 0 5768 400 6 wbs_adr_i[5]
port 34 nsew signal input
rlabel metal2 s 1008 0 1064 400 6 wbs_adr_i[6]
port 35 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 wbs_adr_i[7]
port 36 nsew signal input
rlabel metal2 s 3024 0 3080 400 6 wbs_adr_i[8]
port 37 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 wbs_adr_i[9]
port 38 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 wbs_cyc_i
port 39 nsew signal input
rlabel metal2 s 5376 9600 5432 10000 6 wbs_dat_i[0]
port 40 nsew signal input
rlabel metal3 s 9600 672 10000 728 6 wbs_dat_i[10]
port 41 nsew signal input
rlabel metal3 s 9600 1008 10000 1064 6 wbs_dat_i[11]
port 42 nsew signal input
rlabel metal3 s 9600 1344 10000 1400 6 wbs_dat_i[12]
port 43 nsew signal input
rlabel metal3 s 9600 1680 10000 1736 6 wbs_dat_i[13]
port 44 nsew signal input
rlabel metal3 s 9600 2016 10000 2072 6 wbs_dat_i[14]
port 45 nsew signal input
rlabel metal3 s 9600 2352 10000 2408 6 wbs_dat_i[15]
port 46 nsew signal input
rlabel metal3 s 9600 2688 10000 2744 6 wbs_dat_i[16]
port 47 nsew signal input
rlabel metal3 s 9600 3024 10000 3080 6 wbs_dat_i[17]
port 48 nsew signal input
rlabel metal3 s 9600 3360 10000 3416 6 wbs_dat_i[18]
port 49 nsew signal input
rlabel metal3 s 9600 9744 10000 9800 6 wbs_dat_i[19]
port 50 nsew signal input
rlabel metal3 s 9600 0 10000 56 6 wbs_dat_i[1]
port 51 nsew signal input
rlabel metal3 s 9600 336 10000 392 6 wbs_dat_i[20]
port 52 nsew signal input
rlabel metal3 s 9600 5376 10000 5432 6 wbs_dat_i[21]
port 53 nsew signal input
rlabel metal3 s 9600 5040 10000 5096 6 wbs_dat_i[22]
port 54 nsew signal input
rlabel metal3 s 9600 4704 10000 4760 6 wbs_dat_i[23]
port 55 nsew signal input
rlabel metal3 s 9600 5712 10000 5768 6 wbs_dat_i[24]
port 56 nsew signal input
rlabel metal3 s 9600 6720 10000 6776 6 wbs_dat_i[25]
port 57 nsew signal input
rlabel metal3 s 9600 6384 10000 6440 6 wbs_dat_i[26]
port 58 nsew signal input
rlabel metal3 s 9600 6048 10000 6104 6 wbs_dat_i[27]
port 59 nsew signal input
rlabel metal3 s 9600 7056 10000 7112 6 wbs_dat_i[28]
port 60 nsew signal input
rlabel metal3 s 9600 8064 10000 8120 6 wbs_dat_i[29]
port 61 nsew signal input
rlabel metal3 s 9600 7728 10000 7784 6 wbs_dat_i[2]
port 62 nsew signal input
rlabel metal3 s 9600 7392 10000 7448 6 wbs_dat_i[30]
port 63 nsew signal input
rlabel metal3 s 9600 8400 10000 8456 6 wbs_dat_i[31]
port 64 nsew signal input
rlabel metal3 s 9600 9408 10000 9464 6 wbs_dat_i[3]
port 65 nsew signal input
rlabel metal3 s 9600 9072 10000 9128 6 wbs_dat_i[4]
port 66 nsew signal input
rlabel metal3 s 9600 8736 10000 8792 6 wbs_dat_i[5]
port 67 nsew signal input
rlabel metal2 s 336 9600 392 10000 6 wbs_dat_i[6]
port 68 nsew signal input
rlabel metal2 s 672 9600 728 10000 6 wbs_dat_i[7]
port 69 nsew signal input
rlabel metal2 s 0 9600 56 10000 6 wbs_dat_i[8]
port 70 nsew signal input
rlabel metal2 s 1008 9600 1064 10000 6 wbs_dat_i[9]
port 71 nsew signal input
rlabel metal2 s 2016 9600 2072 10000 6 wbs_dat_o[0]
port 72 nsew signal output
rlabel metal2 s 5712 9600 5768 10000 6 wbs_dat_o[10]
port 73 nsew signal output
rlabel metal2 s 5040 9600 5096 10000 6 wbs_dat_o[11]
port 74 nsew signal output
rlabel metal2 s 6384 9600 6440 10000 6 wbs_dat_o[12]
port 75 nsew signal output
rlabel metal2 s 8064 9600 8120 10000 6 wbs_dat_o[13]
port 76 nsew signal output
rlabel metal2 s 9408 9600 9464 10000 6 wbs_dat_o[14]
port 77 nsew signal output
rlabel metal2 s 9072 9600 9128 10000 6 wbs_dat_o[15]
port 78 nsew signal output
rlabel metal2 s 7392 9600 7448 10000 6 wbs_dat_o[16]
port 79 nsew signal output
rlabel metal2 s 6048 9600 6104 10000 6 wbs_dat_o[17]
port 80 nsew signal output
rlabel metal2 s 1680 9600 1736 10000 6 wbs_dat_o[18]
port 81 nsew signal output
rlabel metal2 s 4704 9600 4760 10000 6 wbs_dat_o[19]
port 82 nsew signal output
rlabel metal2 s 8736 9600 8792 10000 6 wbs_dat_o[1]
port 83 nsew signal output
rlabel metal2 s 7056 9600 7112 10000 6 wbs_dat_o[20]
port 84 nsew signal output
rlabel metal2 s 3360 9600 3416 10000 6 wbs_dat_o[21]
port 85 nsew signal output
rlabel metal2 s 9744 9600 9800 10000 6 wbs_dat_o[22]
port 86 nsew signal output
rlabel metal2 s 8400 9600 8456 10000 6 wbs_dat_o[23]
port 87 nsew signal output
rlabel metal3 s 0 7056 400 7112 6 wbs_dat_o[24]
port 88 nsew signal output
rlabel metal3 s 0 7728 400 7784 6 wbs_dat_o[25]
port 89 nsew signal output
rlabel metal2 s 4032 9600 4088 10000 6 wbs_dat_o[26]
port 90 nsew signal output
rlabel metal2 s 2688 9600 2744 10000 6 wbs_dat_o[27]
port 91 nsew signal output
rlabel metal3 s 0 2688 400 2744 6 wbs_dat_o[28]
port 92 nsew signal output
rlabel metal3 s 0 2352 400 2408 6 wbs_dat_o[29]
port 93 nsew signal output
rlabel metal2 s 6720 9600 6776 10000 6 wbs_dat_o[2]
port 94 nsew signal output
rlabel metal2 s 7728 9600 7784 10000 6 wbs_dat_o[30]
port 95 nsew signal output
rlabel metal2 s 4368 9600 4424 10000 6 wbs_dat_o[31]
port 96 nsew signal output
rlabel metal2 s 3024 9600 3080 10000 6 wbs_dat_o[3]
port 97 nsew signal output
rlabel metal3 s 0 7392 400 7448 6 wbs_dat_o[4]
port 98 nsew signal output
rlabel metal3 s 0 5712 400 5768 6 wbs_dat_o[5]
port 99 nsew signal output
rlabel metal3 s 0 2016 400 2072 6 wbs_dat_o[6]
port 100 nsew signal output
rlabel metal3 s 0 3696 400 3752 6 wbs_dat_o[7]
port 101 nsew signal output
rlabel metal3 s 0 5040 400 5096 6 wbs_dat_o[8]
port 102 nsew signal output
rlabel metal3 s 0 6720 400 6776 6 wbs_dat_o[9]
port 103 nsew signal output
rlabel metal3 s 0 9744 400 9800 6 wbs_sel_i[0]
port 104 nsew signal input
rlabel metal3 s 0 9408 400 9464 6 wbs_sel_i[1]
port 105 nsew signal input
rlabel metal3 s 0 9072 400 9128 6 wbs_sel_i[2]
port 106 nsew signal input
rlabel metal3 s 0 8736 400 8792 6 wbs_sel_i[3]
port 107 nsew signal input
rlabel metal3 s 0 4032 400 4088 6 wbs_stb_i
port 108 nsew signal input
rlabel metal3 s 0 5376 400 5432 6 wbs_we_i
port 109 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 10000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 328002
string GDS_FILE /home/kris/repos/diy-ic/lincoln-gfmpw/openlane/wishbone_register/runs/23_12_05_13_33/results/signoff/wishbone_register.magic.gds
string GDS_START 122518
<< end >>

