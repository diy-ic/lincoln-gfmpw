* NGSPICE file created from titan.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

.subckt titan spi_clock_i spi_cs_i spi_pico_i spi_poci_o sys_clock_i vdd vss
XFILLER_0_27_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7957__A2 _3841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7963_ _1612_ _3841_ _3872_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout56_I net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6914_ _3017_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_53_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7894_ internal_ih.received_byte_count\[5\] internal_ih.received_byte_count\[4\]
+ _3831_ _3834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_119_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6845_ _2953_ ci_adder.uut_simple_neuron.x3\[28\] _2954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8382__A2 _4117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6776_ _2884_ _2885_ _2886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5727_ _1793_ _1834_ _1855_ _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_17_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8515_ ci_adder.output_memory\[12\] _4212_ _4222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8446_ _0704_ _4165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5658_ _1762_ _1788_ _1789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_60_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5589_ _1721_ _1704_ _1717_ _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4609_ _0715_ _0753_ _0772_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8377_ ci_adder.input_memory\[1\]\[6\] _4118_ _4126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7328_ _3357_ _3359_ _3361_ _3362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7259_ ci_adder.uut_simple_neuron.titan_id_1\[3\] ci_adder.uut_simple_neuron.titan_id_0\[3\]
+ _3303_ _3304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7645__A1 ci_adder.uut_simple_neuron.x0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5120__A2 ci_adder.uut_simple_neuron.x2\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__A2 ci_adder.uut_simple_neuron.x3\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8460__I3 _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8373__A2 _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7875__B _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6136__A1 _1960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6611__A2 _2698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4960_ _0909_ _1050_ _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_58_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ _1005_ _1009_ _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6630_ _2738_ _2741_ _2742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8364__A2 _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6561_ _2147_ _2673_ _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_80_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5512_ _1530_ ci_adder.uut_simple_neuron.x2\[30\] _1651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8300_ _3654_ _4071_ _4082_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_119_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6492_ _2252_ _2422_ _2606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6127__A1 _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9305__CLK net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9280_ _0145_ net32 ci_adder.uut_simple_neuron.titan_id_6\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5443_ _1553_ _1583_ _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4689__A1 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8231_ ci_adder.uut_simple_neuron.titan_id_6\[9\] _4046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5374_ _1514_ _1515_ _1516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8162_ ci_adder.output_val_internal\[26\] ci_adder.output_val_internal\[18\] ci_adder.output_val_internal\[10\]
+ ci_adder.output_val_internal\[2\] _3964_ _3961_ _3992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7113_ ci_adder.uut_simple_neuron.titan_id_2\[7\] ci_adder.uut_simple_neuron.titan_id_5\[7\]
+ ci_adder.uut_simple_neuron.titan_id_2\[6\] ci_adder.uut_simple_neuron.titan_id_5\[6\]
+ _3183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__8675__I0 ci_adder.stream_o\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8093_ _3940_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7044_ _3125_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6155__I _2274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8995_ _0478_ net52 spi_interface_cvonk.state\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7946_ _3713_ ci_adder.uut_simple_neuron.x2\[19\] _3855_ _3864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_65_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7695__B ci_adder.uut_simple_neuron.x0\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7877_ internal_ih.instruction_received net13 _3821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_38_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6828_ _2870_ _2937_ _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_92_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8370__I _4116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6759_ _2867_ _2868_ _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8107__A2 _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8429_ _4152_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5341__A2 ci_adder.uut_simple_neuron.x2\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7618__A1 _3599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8291__A1 _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7094__A2 ci_adder.uut_simple_neuron.titan_id_5\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8418__I0 _3746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 ci_adder.uut_simple_neuron.x3\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8280__I _4070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6109__A1 _1807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8656__S _4323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6684__B _2777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5090_ _1217_ _1238_ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8282__A1 ci_adder.uut_simple_neuron.x0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5992_ _2112_ _2114_ _2115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8391__S _4122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8780_ _0327_ net25 ci_adder.uut_simple_neuron.x2\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_7800_ _3754_ _3755_ _3756_ _3757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_93_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4943_ _1055_ _1091_ _1092_ _1095_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_7731_ _3524_ _3695_ _3699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_86_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7662_ ci_adder.uut_simple_neuron.x3\[5\] _3617_ _3642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6613_ _2677_ _2687_ _2724_ _2725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4874_ _1027_ _1028_ _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout19_I net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7593_ ci_adder.uut_simple_neuron.x0\[27\] ci_adder.uut_simple_neuron.x0\[28\] _3581_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6544_ _2471_ _2657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6475_ _2548_ _2550_ _2589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7699__I1 ci_adder.uut_simple_neuron.x3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9263_ _0158_ net64 ci_adder.uut_simple_neuron.titan_id_6\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5426_ _1484_ _1486_ _1533_ _1567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8214_ _4037_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6520__A1 _1723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8845__CLK net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9194_ _0088_ net64 ci_adder.uut_simple_neuron.titan_id_2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5357_ _0993_ _1499_ _1500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8145_ _3824_ _3976_ _3977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5288_ _1409_ _1413_ _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8076_ internal_ih.byte6\[1\] internal_ih.byte5\[1\] _3930_ _3932_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5626__A3 _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7027_ _3110_ _3111_ _3112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8995__CLK net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6587__A1 _2648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8978_ _0461_ net35 ci_adder.uut_simple_neuron.x0\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7929_ _3840_ _3855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_93_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8328__A2 _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6339__A1 _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5011__A1 ci_adder.uut_simple_neuron.x2\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8500__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8639__I0 ci_adder.stream_o\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5078__A1 ci_adder.uut_simple_neuron.x2\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9000__CLK net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9150__CLK net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5250__A1 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5002__A1 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5553__A2 _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4590_ _0744_ _0746_ _0754_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_25_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8868__CLK net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6260_ _2276_ _2313_ _2377_ _2378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_40_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6191_ _2296_ _2309_ _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_86_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5211_ _1233_ ci_adder.uut_simple_neuron.x2\[22\] _1354_ _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5142_ _1285_ _1289_ _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5069__A1 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5073_ _0712_ _1221_ _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8901_ _0060_ net13 ci_adder.value_i\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_48_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8832_ _0379_ net21 internal_ih.byte6\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5241__A1 _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ ci_adder.uut_simple_neuron.x3\[16\] _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8763_ _0310_ net81 ci_adder.uut_simple_neuron.x2\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4926_ _0908_ _1050_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7714_ _3619_ _3683_ _3684_ _3685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8694_ _4346_ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4857_ _0874_ _0974_ _1006_ _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_47_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7645_ ci_adder.uut_simple_neuron.x0\[3\] _3623_ _3627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_118_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7576_ _3567_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6527_ _2523_ _2569_ _2641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6741__A1 _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4788_ _0925_ _0944_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_15_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9315_ _0576_ net22 ci_adder.stream_o\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6458_ _2451_ _2500_ _2573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9246_ _0111_ net78 ci_adder.uut_simple_neuron.titan_id_5\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9177_ _0210_ net79 ci_adder.uut_simple_neuron.titan_id_3\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6389_ _2389_ _2441_ _2505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5409_ _0994_ _1543_ _1550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9023__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8128_ _3811_ _3960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__9173__CLK net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8059_ internal_ih.byte5\[1\] internal_ih.byte4\[1\] _3919_ _3923_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8021__I1 internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8572__I2 ci_adder.uut_simple_neuron.x2\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9041__D ci_adder.input_memory\[1\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5760_ _1883_ _1887_ _1888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5691_ _1816_ _1820_ _1821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4711_ _0845_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_57_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4642_ _0710_ _0790_ _0785_ _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7430_ ci_adder.uut_simple_neuron.titan_id_1\[2\] ci_adder.uut_simple_neuron.titan_id_0\[2\]
+ _3446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4573_ _0710_ _0724_ _0734_ _0735_ _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_7361_ ci_adder.uut_simple_neuron.titan_id_1\[19\] ci_adder.uut_simple_neuron.titan_id_0\[19\]
+ _3389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9046__CLK net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6312_ _2420_ _2426_ _2428_ _2429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7292_ _3331_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9100_ _0195_ net64 ci_adder.uut_simple_neuron.titan_id_0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout7 net11 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8476__A1 _4165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6243_ _2300_ _2360_ _2361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_12_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9031_ _0514_ net43 internal_ih.expected_byte_count\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6174_ _1882_ _2292_ _2293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout86_I net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5125_ _1263_ _1266_ _1272_ _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5056_ _1203_ _1172_ _1205_ _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7451__A2 _3459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_88_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8815_ _0362_ net23 internal_ih.byte4\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5958_ _1723_ _1757_ _2081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8746_ _0293_ net44 internal_ih.received_byte_count\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4909_ _1036_ _1062_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5889_ _1976_ _1975_ _2014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_90_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8554__I2 ci_adder.uut_simple_neuron.x2\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8677_ ci_adder.stream_o\[23\] ci_adder.output_memory\[23\] _4334_ _4338_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6714__A1 _2364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7628_ _3599_ _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7559_ _3547_ _3550_ _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9229_ _0123_ net86 ci_adder.uut_simple_neuron.titan_id_5\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8562__S1 _4253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7722__I _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8553__I _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9069__CLK net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7632__I _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8906__CLK net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8664__S _4323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5444__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6930_ _3010_ _3019_ _3030_ _3031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6861_ _0163_ _2930_ _2970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5812_ _1902_ _1938_ _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6792_ _2304_ _2901_ _2902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8600_ _4257_ _4288_ _4290_ _4291_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__5747__A2 _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5743_ _1702_ _1752_ _1870_ _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_85_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8531_ ci_adder.uut_simple_neuron.x0\[15\] ci_adder.input_memory\[1\]\[15\] _1011_
+ _2050_ _4206_ _4207_ _4235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_57_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8536__I2 ci_adder.uut_simple_neuron.x2\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5674_ ci_adder.uut_simple_neuron.x3\[8\] ci_adder.uut_simple_neuron.x3\[9\] _1804_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8462_ ci_adder.output_val_internal\[2\] _4170_ _4179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4625_ ci_adder.uut_simple_neuron.x2\[6\] _0787_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7413_ _3427_ _3428_ _3431_ _3432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8393_ _3685_ ci_adder.input_memory\[1\]\[14\] _4122_ _4134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4556_ _0710_ _0715_ _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7344_ _3371_ _3372_ _3374_ _3375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7275_ ci_adder.uut_simple_neuron.titan_id_1\[6\] ci_adder.uut_simple_neuron.titan_id_0\[6\]
+ _3317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4487_ _0597_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6226_ _2342_ _2343_ _2344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9014_ _0497_ net36 ci_adder.input_memory\[1\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7672__A2 _3619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6157_ _2228_ _2234_ _2275_ _2276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5108_ _1252_ _1254_ _1255_ _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__8621__A1 _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5997__I _2119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6088_ _2205_ _2208_ _2209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5039_ _1182_ _1188_ _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_28_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9211__CLK net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8480__S0 _4166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7983__I0 internal_ih.byte0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8729_ spi_interface_cvonk.SCLK_r\[1\] net44 spi_interface_cvonk.SCLK_r\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8929__CLK net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8548__I _4161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7663__A2 _3641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5674__A1 ci_adder.uut_simple_neuron.x3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4477__A2 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7627__I _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4401__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4410_ _0629_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_124_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5390_ _0711_ _1531_ _1532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__S1 _4207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7060_ ci_adder.uut_simple_neuron.titan_id_4\[30\] ci_adder.uut_simple_neuron.titan_id_3\[30\]
+ _3139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7654__A2 _3608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6011_ _2089_ _2131_ _2132_ _2133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9234__CLK net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5417__A1 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7962_ _3751_ _3846_ _3872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6913_ _3015_ _3016_ _3017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout49_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7893_ internal_ih.received_byte_count\[4\] _3831_ internal_ih.received_byte_count\[5\]
+ _3833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6844_ ci_adder.uut_simple_neuron.x3\[27\] _2953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6775_ _2817_ _2821_ _2885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5726_ _1837_ _1854_ _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8514_ _4211_ _4218_ _4220_ _4221_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_94_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8445_ ci_adder.output_memory\[0\] _4163_ _4164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5657_ _1785_ _1787_ _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_72_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5588_ _1699_ _1721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_96_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4608_ _0709_ _0766_ _0768_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8376_ _3641_ _4117_ _4125_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7327_ ci_adder.uut_simple_neuron.titan_id_1\[13\] ci_adder.uut_simple_neuron.titan_id_0\[13\]
+ _3361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4539_ _0689_ _0701_ _0708_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_68_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8693__I1 ci_adder.output_memory\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7258_ ci_adder.uut_simple_neuron.titan_id_1\[2\] ci_adder.uut_simple_neuron.titan_id_0\[2\]
+ _3303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6209_ _2323_ _2324_ _2325_ _2327_ _2328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_7189_ ci_adder.uut_simple_neuron.titan_id_2\[21\] ci_adder.uut_simple_neuron.titan_id_5\[21\]
+ _3246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_5_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__A1 _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6351__I ci_adder.uut_simple_neuron.x3\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7708__I0 ci_adder.value_i\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9107__CLK net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7884__A2 _3826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_39_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7636__A2 _3599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4890_ _1041_ _1018_ _1043_ _0976_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_73_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6560_ _2249_ _2607_ _2606_ _2673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_80_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5511_ _1530_ ci_adder.uut_simple_neuron.x2\[30\] _1650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6491_ _2252_ _2422_ _2605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8389__S _4122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5442_ _1470_ _1582_ _1583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_57_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8230_ _4045_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5373_ _1470_ _1497_ _1515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8161_ _3963_ ci_adder.stream_o\[2\] ci_adder.stream_o\[18\] _3965_ _3990_ _3991_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__9224__D _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7112_ _3180_ _3181_ _3182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8092_ internal_ih.byte7\[1\] internal_ih.byte6\[1\] _3930_ _3940_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7043_ _3122_ _3124_ _3125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_2_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_66_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8994_ _0477_ net52 spi_interface_cvonk.state\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7945_ _1161_ _3841_ _3863_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7938__I0 _3691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7876_ _3811_ _3819_ _3820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_6827_ _2874_ _2936_ _2937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_65_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6758_ _2792_ _2865_ _2868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6689_ _2728_ _2753_ _2800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5709_ _1801_ _1807_ _1838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8428_ _3768_ ci_adder.input_memory\[1\]\[31\] _4116_ _4152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8359_ _3781_ _4109_ spi_interface_cvonk.state\[2\] _4115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5341__A3 ci_adder.uut_simple_neuron.x2\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7618__A2 _3601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8291__A2 _4072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8561__I _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6357__A2 _2423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7905__I _3840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7857__A2 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8282__A2 _4072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6293__A1 _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8797__CLK net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5991_ _2026_ _2063_ _2113_ _2114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_78_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4942_ _1093_ _1094_ _1089_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7730_ _3698_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7661_ ci_adder.value_i\[5\] _3619_ _3640_ _3641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6612_ _2654_ _2676_ _2724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4873_ _0992_ _0995_ _1026_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7545__A1 _3524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4359__A1 internal_ih.current_instruction\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7592_ _3580_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6543_ _2604_ _2608_ _2655_ _2656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6474_ _2557_ _2567_ _2587_ _2588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9262_ _0157_ net64 ci_adder.uut_simple_neuron.titan_id_6\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5425_ _0712_ ci_adder.uut_simple_neuron.x2\[27\] _1530_ _1566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8213_ ci_adder.uut_simple_neuron.titan_id_6\[0\] _4037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9193_ _0077_ net63 ci_adder.uut_simple_neuron.titan_id_2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5356_ _1467_ _1498_ _1499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8144_ internal_ih.spi_rx_byte_i\[2\] _3806_ _3976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5287_ _1397_ _1408_ _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8075_ _3931_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7026_ ci_adder.uut_simple_neuron.titan_id_4\[25\] ci_adder.uut_simple_neuron.titan_id_3\[25\]
+ _3111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XPHY_EDGE_ROW_74_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8977_ _0460_ net35 ci_adder.uut_simple_neuron.x0\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7928_ _3667_ _3842_ _3854_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6339__A2 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9129__D _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7859_ _3801_ _3803_ _3775_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_108_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_83_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5011__A2 ci_adder.uut_simple_neuron.x2\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8336__I0 _3746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8639__I1 ci_adder.output_memory\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6027__A1 _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7635__I _3608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5210_ _1351_ _1355_ _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6190_ _2305_ _2308_ _2309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5141_ _1207_ _1286_ _1288_ _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5072_ _1220_ _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8900_ _0059_ net13 ci_adder.value_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7766__A1 _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8831_ _0378_ net21 internal_ih.byte6\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8762_ _0309_ net81 ci_adder.uut_simple_neuron.x2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5974_ ci_adder.uut_simple_neuron.x3\[13\] _2095_ _2096_ _2097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA_fanout31_I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7713_ ci_adder.value_i\[14\] _3659_ _3684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4925_ _1054_ _1060_ _1077_ _1042_ _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_59_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8693_ ci_adder.stream_o\[31\] ci_adder.output_memory\[31\] _3601_ _4346_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4856_ ci_adder.uut_simple_neuron.x2\[15\] _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7644_ _3612_ _3625_ _3626_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8812__CLK net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7575_ _3563_ _3566_ _3567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8318__I0 _3703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6526_ _2583_ _2586_ _2639_ _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_4787_ _0927_ _0930_ _0943_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_16_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9314_ _0575_ net45 ci_adder.stream_o\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6457_ _2451_ _2500_ _2572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9245_ _0110_ net78 ci_adder.uut_simple_neuron.titan_id_5\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_31_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8962__CLK net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6388_ _2501_ _2503_ _2504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_100_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5408_ _1516_ _1542_ _1549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9176_ _0209_ net75 ci_adder.uut_simple_neuron.titan_id_3\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5339_ _1480_ _1481_ _1482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_8127_ _3815_ _3959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__9318__CLK net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8058_ _3922_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7009_ _3096_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8572__I3 _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6248__A1 ci_adder.uut_simple_neuron.x3\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6799__A2 _2825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8835__CLK net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5690_ _1817_ _1818_ _1819_ _1820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4982__A1 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4710_ _0847_ _0858_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4641_ _0753_ _0770_ _0802_ _0795_ _0786_ _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7920__A1 _3645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4734__B2 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4572_ _0737_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7360_ _3381_ _3386_ _3388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_13_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6311_ _2097_ _2427_ _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7291_ _3329_ _3330_ _3331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8397__S _4122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout8 net11 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6242_ _2200_ _2301_ _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6487__A1 _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9030_ _0513_ net43 internal_ih.expected_byte_count\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6239__A1 _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6173_ _1958_ _2256_ _2291_ _2292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_fanout79_I net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5124_ _1270_ _1271_ _1272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5055_ _1174_ _1204_ _1205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_88_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8814_ _0361_ net16 internal_ih.byte3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5957_ _1723_ _1757_ _2080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_94_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8745_ _0292_ net43 internal_ih.received_byte_count\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4908_ _1040_ _1044_ _1061_ _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__4973__A1 _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8676_ _4337_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5888_ _2012_ _1974_ _2013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7627_ _3611_ _3612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8554__I3 _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4839_ _0993_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7911__A1 _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7208__C ci_adder.uut_simple_neuron.titan_id_5\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7558_ ci_adder.uut_simple_neuron.x0\[21\] ci_adder.uut_simple_neuron.x0\[22\] _3552_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6509_ _2087_ _2105_ _2623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7489_ _3488_ _3491_ _3494_ _3495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8467__A2 _4170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9140__CLK net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9228_ _0122_ net85 ci_adder.uut_simple_neuron.titan_id_5\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8100__S _3825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5150__A1 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9142__D _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9159_ _0159_ net66 ci_adder.uut_simple_neuron.titan_id_3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9290__CLK net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6650__A1 _1807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8490__I2 ci_adder.uut_simple_neuron.x2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8858__CLK net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Left_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4964__A1 _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6860_ _2927_ _2929_ _2969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5811_ _1903_ _1937_ _1938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6791_ _2422_ _2820_ _2819_ _2901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9013__CLK net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5742_ _1849_ _1850_ _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7992__I1 internal_ih.byte0\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8530_ ci_adder.output_memory\[15\] _4212_ _4234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5673_ ci_adder.uut_simple_neuron.x3\[6\] _1775_ _1802_ _1803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_60_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8536__I3 _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8461_ _4165_ _4177_ _4178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8392_ _4133_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4624_ ci_adder.uut_simple_neuron.x2\[7\] _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7412_ _3430_ _3431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4555_ ci_adder.uut_simple_neuron.x2\[3\] _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7343_ ci_adder.uut_simple_neuron.titan_id_1\[16\] ci_adder.uut_simple_neuron.titan_id_0\[16\]
+ _3374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9013_ _0496_ net37 ci_adder.input_memory\[1\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7274_ _3313_ _3315_ _3316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4486_ _0669_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6225_ _0163_ _2285_ _2343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6156_ _2231_ _2233_ _2275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5107_ _1223_ _1253_ _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6087_ _2207_ _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5038_ _1186_ _1187_ _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_28_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5199__A1 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6989_ ci_adder.uut_simple_neuron.titan_id_4\[16\] ci_adder.uut_simple_neuron.titan_id_3\[16\]
+ _3080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8480__S1 _4167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8728_ spi_interface_cvonk.SCLK_r\[0\] net43 spi_interface_cvonk.SCLK_r\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7934__S _3855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8659_ _4328_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6699__A1 ci_adder.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5123__A1 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5674__A2 ci_adder.uut_simple_neuron.x3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6623__A1 ci_adder.uut_simple_neuron.x3\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9036__CLK net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8376__A1 _3641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4937__A1 _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7103__A2 ci_adder.uut_simple_neuron.titan_id_5\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8300__A1 _3654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5114__A1 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6010_ _2092_ _2107_ _2132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input3_I spi_pico_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8603__A2 _4293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7961_ _1485_ _3841_ _3871_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_85_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5112__B _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6912_ ci_adder.uut_simple_neuron.titan_id_4\[6\] ci_adder.uut_simple_neuron.titan_id_3\[6\]
+ _3016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7892_ _3826_ _3832_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6843_ _2950_ _2951_ _2952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8367__A1 _3621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6774_ _2808_ _2816_ _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4928__A1 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5725_ _1839_ _1853_ _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_73_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout8_I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8513_ ci_adder.output_val_internal\[11\] _4203_ _4221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5656_ _1722_ _1763_ _1743_ _1786_ _1787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_45_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8444_ _0703_ _4163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_115_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4607_ _0715_ _0742_ _0753_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_5_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8649__I _3601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5587_ _1720_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_96_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8375_ ci_adder.input_memory\[1\]\[5\] _4118_ _4125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7326_ _3360_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4538_ _0689_ _0707_ ci_adder.stream_enabled _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4469_ internal_ih.byte1\[3\] _0659_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7257_ _3302_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6208_ _2271_ _2326_ _2327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6853__A1 ci_adder.uut_simple_neuron.x3\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7188_ _3243_ _3244_ _3245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9059__CLK net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6139_ _2255_ _2258_ _2259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_84_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5592__A1 _1723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8125__A4 _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8559__I _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6072__A2 _2147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_103_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4622__A3 ci_adder.uut_simple_neuron.x2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5583__A1 _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5510_ _1647_ _1625_ _1648_ _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6490_ _2596_ _2603_ _2604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_81_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5441_ _1556_ _1581_ _1582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5335__A1 ci_adder.uut_simple_neuron.x2\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5372_ _1473_ _1496_ _1514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8160_ _3966_ _3989_ _3990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7111_ _3170_ _3174_ _3181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8091_ _3939_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7042_ _3119_ _3120_ _3123_ _3124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5638__A2 _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout61_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8993_ _0476_ net45 internal_ih.data_pointer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7944_ _3708_ _3846_ _3863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8919__CLK net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7938__I1 _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7875_ internal_ih.instruction_received _3816_ _3818_ _3819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6826_ _2876_ _2935_ _2936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_65_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6757_ _2794_ _2864_ _2867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5574__A1 _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5708_ _1677_ _1836_ _1837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_98_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6688_ _2766_ _2779_ _2798_ _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5639_ _1686_ _1769_ _1770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5326__A1 _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8427_ _4151_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8358_ _3780_ _3782_ _4114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7309_ _3344_ _3345_ _3346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8289_ _3631_ _4076_ _4077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5565__A1 _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9224__CLK net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5990_ _2029_ _2062_ _2113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4941_ ci_adder.uut_simple_neuron.x2\[15\] ci_adder.uut_simple_neuron.x2\[16\] ci_adder.uut_simple_neuron.x2\[17\]
+ _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_47_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4872_ _0992_ _0995_ _1026_ _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_24_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7660_ _3608_ _3638_ _3639_ _3640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6611_ _2721_ _2698_ _2722_ _2723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7591_ _3576_ _3579_ _3580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6542_ _2596_ _2603_ _2655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6473_ _2533_ _2556_ _2587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9261_ _0156_ net64 ci_adder.uut_simple_neuron.titan_id_6\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5424_ _1482_ _1563_ _1564_ _1487_ _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_8212_ _3979_ _4035_ _4036_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9192_ _0066_ net50 ci_adder.uut_simple_neuron.titan_id_2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8143_ internal_ih.spi_rx_byte_i\[1\] _3812_ _3974_ _3975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5355_ _1470_ _1497_ _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5286_ _1119_ _1428_ _1429_ _1430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8074_ internal_ih.byte6\[0\] internal_ih.byte5\[0\] _3930_ _3931_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7025_ ci_adder.uut_simple_neuron.titan_id_4\[24\] ci_adder.uut_simple_neuron.titan_id_3\[24\]
+ _3099_ _3107_ _3109_ _3110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__7481__A1 ci_adder.uut_simple_neuron.x0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8741__CLK net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8976_ _0459_ net37 ci_adder.uut_simple_neuron.x0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5795__A1 _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7927_ ci_adder.uut_simple_neuron.x2\[10\] _3846_ _3854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7858_ spi_interface_cvonk.buffer\[7\] _3802_ _3776_ _3803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6809_ _2850_ _2852_ _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7789_ _3747_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7942__S _3855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8592__S0 _4252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4586__B ci_adder.uut_simple_neuron.x2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6027__A2 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8013__S _3897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ _1246_ _1287_ _1244_ _1288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5071_ _1161_ _1184_ _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7463__A1 _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6018__A2 _2100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8830_ _0377_ net15 internal_ih.byte5\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5777__A1 _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5973_ ci_adder.uut_simple_neuron.x3\[14\] _2050_ _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7766__A2 _3632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8761_ _0308_ net81 ci_adder.uut_simple_neuron.x2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_48_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4924_ _0714_ _1058_ _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7712_ _3508_ _3682_ _3683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8015__I0 internal_ih.byte2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8692_ _4345_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ _0808_ _1005_ _1009_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7643_ _1679_ _3617_ _3626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout24_I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4786_ _0934_ _0942_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7574_ _3564_ _3565_ _3566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6525_ _2628_ _2638_ _2639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4752__A2 _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9313_ _0574_ net22 ci_adder.stream_o\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8318__I1 _3524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9244_ _0109_ net79 ci_adder.uut_simple_neuron.titan_id_5\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_16_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ _2520_ _2570_ _2571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6387_ _2391_ _2440_ _2502_ _2503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5407_ _1548_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9175_ _0208_ net90 ci_adder.uut_simple_neuron.titan_id_3\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5338_ _1221_ _1352_ _1398_ _1481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_8126_ _3957_ _3958_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7454__A1 _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8057_ internal_ih.byte5\[0\] internal_ih.byte4\[0\] _3919_ _3922_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7008_ ci_adder.uut_simple_neuron.titan_id_4\[22\] ci_adder.uut_simple_neuron.titan_id_3\[22\]
+ _3095_ _3096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5269_ _1409_ _1413_ _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8959_ _0032_ net7 ci_adder.instruction_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8006__I0 internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7693__A1 ci_adder.uut_simple_neuron.x3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6248__A2 _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4431__B2 internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4640_ _0792_ _0793_ _0713_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_72_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7920__A2 _3841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6310_ _2100_ _2249_ _2427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4571_ _0734_ _0736_ _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_52_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7290_ ci_adder.uut_simple_neuron.titan_id_1\[8\] ci_adder.uut_simple_neuron.titan_id_0\[8\]
+ _3330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout9 net11 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6241_ _2305_ _2308_ _2358_ _2359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_90_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6172_ _1960_ _2097_ _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4498__A1 internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6239__A2 _2356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5123_ _0712_ _1234_ _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5054_ _1145_ _1202_ _1172_ _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_88_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8813_ _0360_ net18 internal_ih.byte3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5956_ _2077_ _2078_ _2079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8744_ _0291_ net43 internal_ih.received_byte_count\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5887_ _1971_ _2012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4907_ _1054_ _1060_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8675_ ci_adder.stream_o\[22\] ci_adder.output_memory\[22\] _4334_ _4337_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6175__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4838_ _0870_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_23_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7626_ _3607_ _3610_ _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_35_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7911__A2 _3841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5922__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ _0808_ _0852_ _0910_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7557_ _3551_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_120_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6508_ _2620_ _2554_ _2621_ _2622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7488_ ci_adder.uut_simple_neuron.x0\[9\] ci_adder.uut_simple_neuron.x0\[10\] _3494_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6439_ _2053_ _2553_ _2554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9227_ _0121_ net85 ci_adder.uut_simple_neuron.titan_id_5\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7675__A1 _3479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9158_ ci_adder.uut_simple_neuron.x2\[0\] net48 ci_adder.uut_simple_neuron.titan_id_3\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8109_ internal_ih.spi_rx_byte_i\[1\] internal_ih.current_instruction\[1\] _3947_
+ _3949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8475__I0 _3459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9089_ _0542_ net34 ci_adder.output_val_internal\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8490__I3 ci_adder.uut_simple_neuron.x3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6166__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6469__A2 _2527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7666__A1 ci_adder.value_i\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_72_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8802__CLK net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4652__A1 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5810_ _1933_ _1936_ _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6790_ _2899_ _2900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8952__CLK net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5741_ _1837_ _1854_ _1868_ _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_57_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8460_ ci_adder.uut_simple_neuron.x0\[2\] ci_adder.input_memory\[1\]\[2\] _0724_
+ _1679_ _4166_ _4167_ _4177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_45_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5672_ ci_adder.uut_simple_neuron.x3\[7\] ci_adder.uut_simple_neuron.x3\[8\] _1802_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7411_ ci_adder.uut_simple_neuron.titan_id_1\[28\] ci_adder.uut_simple_neuron.titan_id_0\[28\]
+ _3430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9308__CLK net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4623_ _0784_ _0785_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_72_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8391_ _3680_ ci_adder.input_memory\[1\]\[13\] _4122_ _4133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7342_ _3373_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4554_ _0721_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7657__A1 _3612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7273_ _3311_ _3314_ _3315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout91_I net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6224_ _1871_ _1886_ _2342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9012_ _0495_ net37 ci_adder.input_memory\[1\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4485_ internal_ih.byte2\[3\] _0659_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_0_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6155_ _2274_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6086_ _1917_ _2206_ _2207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5106_ _1223_ _1253_ _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5037_ _1159_ _1162_ _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_68_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8385__A2 _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8670__I _3601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6988_ _3071_ _3076_ _3079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8727_ net1 net43 spi_interface_cvonk.SCLK_r\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5939_ _2029_ _2062_ _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6404__B _2457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8658_ ci_adder.stream_o\[14\] ci_adder.output_memory\[14\] _4323_ _4328_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7609_ _3594_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8589_ ci_adder.output_val_internal\[25\] _4249_ _4283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7648__A1 ci_adder.value_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7950__S _3855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8825__CLK net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6623__A2 ci_adder.uut_simple_neuron.x3\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8975__CLK net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6387__A1 _2391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8376__A2 _4117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4937__A2 ci_adder.uut_simple_neuron.x2\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7887__A1 _3826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8021__S _3897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7639__A1 _3612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8300__A2 _4071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7960_ _3746_ _3846_ _3871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8691__S _3601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6911_ _3013_ _3014_ _3015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7891_ internal_ih.received_byte_count\[4\] _3831_ _3832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6842_ _2896_ _2897_ _2951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8367__A2 _4117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9130__CLK net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6773_ _2824_ _2827_ _2882_ _2883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8119__A2 _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5724_ _1848_ _1852_ _1853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8512_ _4214_ _4219_ _4220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5655_ _1759_ _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8443_ _4161_ _4162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4606_ _0766_ _0769_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_8374_ _3636_ _4117_ _4124_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6550__A1 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5586_ _1717_ _1719_ _1720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7325_ _3357_ _3359_ _3360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8848__CLK net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4537_ _0704_ _0706_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6302__A1 _2364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4468_ _0660_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7256_ ci_adder.uut_simple_neuron.titan_id_2\[0\] ci_adder.uut_simple_neuron.titan_id_5\[0\]
+ _3302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6207_ _2272_ _2326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6853__A2 _2356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7187_ _3240_ _3241_ _3244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6138_ _2257_ _2258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_5_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4399_ internal_ih.byte4\[2\] _0623_ _0620_ internal_ih.byte0\[2\] _0624_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_99_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6069_ _1878_ _2149_ _2189_ _2190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_95_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8530__A2 _4212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8294__A1 _3641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4855__A1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9153__CLK net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4607__A1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4622__A4 ci_adder.uut_simple_neuron.x2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5032__A1 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6780__A1 ci_adder.uut_simple_neuron.x3\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5440_ _1560_ _1580_ _1581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5371_ _1422_ _1508_ _1509_ _1512_ _1513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8090_ internal_ih.byte7\[0\] internal_ih.byte6\[0\] _3930_ _3939_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8285__A1 _3621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7110_ _3178_ _3179_ _3168_ _3180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7041_ ci_adder.uut_simple_neuron.titan_id_4\[27\] ci_adder.uut_simple_neuron.titan_id_3\[27\]
+ _3123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8992_ _0475_ net18 ci_adder.uut_simple_neuron.x0\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8588__A2 _4281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7943_ _3862_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout54_I net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7874_ _3817_ _3782_ _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_9_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6825_ _2879_ _2934_ _2935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6756_ _2866_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5574__A2 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5707_ _1692_ _1730_ _1835_ _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_98_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6687_ _2725_ _2765_ _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5638_ _1681_ _1711_ _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8426_ _3765_ ci_adder.input_memory\[1\]\[30\] _4116_ _4151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5569_ _1677_ _1703_ _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_60_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8357_ _4111_ _3781_ _4112_ _4109_ _4113_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__9026__CLK net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7308_ _3341_ _3342_ _3345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8288_ _4070_ _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__9176__CLK net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7239_ ci_adder.uut_simple_neuron.titan_id_2\[28\] ci_adder.uut_simple_neuron.titan_id_5\[28\]
+ _3288_ _3289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_87_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5014__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4828__A1 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5253__A1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4940_ _1011_ ci_adder.uut_simple_neuron.x2\[16\] _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_35_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4871_ _0996_ _1025_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5005__A1 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8042__I1 internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6610_ _2652_ _2688_ _2722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_74_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7590_ _3573_ _3577_ _3578_ _3572_ _3579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_15_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6541_ _2610_ _2614_ _2653_ _2654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9049__CLK net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6472_ _2528_ _2584_ _2585_ _2586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_54_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9260_ _0155_ net63 ci_adder.uut_simple_neuron.titan_id_6\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5423_ _1530_ _1488_ _1564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8211_ internal_ih.spi_tx_byte_o\[7\] _3978_ _4036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9191_ ci_adder.uut_simple_neuron.titan_id_0\[1\] net49 ci_adder.uut_simple_neuron.titan_id_2\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5354_ _1473_ _1496_ _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9199__CLK net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8142_ internal_ih.instruction_received _0599_ _3819_ _3974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_10_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5285_ _1084_ _1412_ _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9251__D _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8073_ _3818_ _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7024_ _3108_ _3109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8975_ _0458_ net60 ci_adder.uut_simple_neuron.x0\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5795__A2 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7926_ _3853_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7857_ _3786_ _3784_ _3802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6808_ _2881_ _2917_ _2918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_122_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7788_ _3746_ ci_adder.uut_simple_neuron.x3\[26\] _3692_ _3747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _2848_ _2849_ _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8592__S1 _4253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8409_ _4142_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout90 net91 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_83_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8909__CLK net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5070_ _0808_ _1083_ _1218_ _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7463__A2 _3470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5777__A2 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5972_ ci_adder.uut_simple_neuron.x3\[14\] _2050_ _2095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8760_ _0307_ net58 ci_adder.uut_simple_neuron.x2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_48_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4923_ _1047_ _1053_ _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7711_ ci_adder.uut_simple_neuron.x0\[12\] _3502_ _3670_ _3682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__8015__I1 internal_ih.byte1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8691_ ci_adder.stream_o\[30\] ci_adder.output_memory\[30\] _3601_ _4345_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4854_ _0939_ _1008_ _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7642_ ci_adder.value_i\[2\] _3613_ _3624_ _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4785_ _0935_ _0926_ _0941_ _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_7573_ _3556_ _3559_ _3565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout17_I net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6524_ _2629_ _2637_ _2638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9312_ _0573_ net22 ci_adder.stream_o\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8479__A1 ci_adder.output_memory\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9243_ _0108_ net79 ci_adder.uut_simple_neuron.titan_id_5\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_70_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6455_ _2523_ _2569_ _2570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_31_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6386_ _2394_ _2439_ _2502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5406_ _1513_ _1547_ _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9174_ _0207_ net90 ci_adder.uut_simple_neuron.titan_id_3\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5337_ _1447_ _1479_ _1480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8125_ _3807_ _3808_ _3814_ _3818_ _3958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5268_ _1084_ _1151_ _1412_ _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7454__A2 _3459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8056_ _3921_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7007_ _3091_ _3092_ _3094_ _3095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_76_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5199_ _0714_ _1270_ _1345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9214__CLK net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8958_ _0031_ net7 ci_adder.instruction_i\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7909_ _3621_ _3841_ _3844_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8889_ _0436_ net33 ci_adder.output_memory\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5537__I ci_adder.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7693__A2 _3632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5208__A1 ci_adder.uut_simple_neuron.x2\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4431__A2 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4570_ _0710_ _0724_ _0735_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8731__CLK net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5931__A2 _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6240_ _2298_ _2304_ _2358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7684__A2 _3659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5182__I _1328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6171_ _2242_ _2260_ _2289_ _2290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_90_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5122_ _1221_ _1267_ _1269_ _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_20_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5053_ _1145_ _1202_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_88_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8812_ _0359_ net17 internal_ih.byte3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5955_ _1728_ _2041_ _2078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8743_ _0290_ net44 spi_interface_cvonk.buffer\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5886_ _2008_ _2010_ _2011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_117_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4906_ _1059_ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8674_ _4336_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4837_ _0953_ _0982_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7625_ _3608_ _3609_ _3610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5922__A2 _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4768_ _0923_ _0924_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7556_ _3547_ _3550_ _3551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6507_ _2090_ _2553_ _2621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4699_ _0847_ _0858_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7487_ ci_adder.uut_simple_neuron.x0\[11\] _3493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_15_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6438_ _2143_ _2480_ _2552_ _2553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9226_ _0120_ net85 ci_adder.uut_simple_neuron.titan_id_5\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9157_ _0249_ net76 ci_adder.uut_simple_neuron.titan_id_4\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6369_ _2097_ _2427_ _2484_ _2485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8108_ _0596_ _3947_ _3948_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9088_ _0541_ net34 ci_adder.output_val_internal\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8109__S _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8039_ _3912_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7948__S _3855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4413__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7666__A2 _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5429__A1 ci_adder.uut_simple_neuron.x2\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8615__A1 _4170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8019__S _3897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4652__A2 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5740_ _1839_ _1853_ _1868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7729__I0 _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5671_ _1713_ _1777_ _1800_ _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7410_ _3429_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_20_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4622_ ci_adder.uut_simple_neuron.x2\[2\] ci_adder.uut_simple_neuron.x2\[3\] ci_adder.uut_simple_neuron.x2\[4\]
+ ci_adder.uut_simple_neuron.x2\[5\] _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_8390_ _4132_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4553_ _0719_ _0720_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7341_ _3371_ _3372_ _3373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_52_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7657__A2 _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7272_ ci_adder.uut_simple_neuron.titan_id_1\[5\] ci_adder.uut_simple_neuron.titan_id_0\[5\]
+ _3314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_4_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4484_ _0668_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5668__A1 _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6223_ _2288_ _2339_ _2340_ _2341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9011_ _0494_ net37 ci_adder.input_memory\[1\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6154_ _2271_ _2273_ _2274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout84_I net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8437__B _3966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8606__A1 ci_adder.output_memory\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6085_ _1919_ _2049_ _2206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5105_ _1232_ _1236_ _1253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5036_ _1183_ _1185_ _1186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8777__CLK net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_28_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8465__S0 _4166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6987_ ci_adder.uut_simple_neuron.titan_id_4\[18\] ci_adder.uut_simple_neuron.titan_id_3\[18\]
+ _3078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_0_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5938_ _2035_ _2061_ _2062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8726_ _0281_ net18 ci_adder.uut_simple_neuron.x3\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5869_ _1958_ _1960_ _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_106_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8657_ _4327_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7608_ _3592_ _3593_ _3594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8588_ _4260_ _4281_ _4282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7539_ _3524_ ci_adder.uut_simple_neuron.x0\[18\] _3532_ _3537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_114_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7648__A2 _3629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9209_ _0074_ net74 ci_adder.uut_simple_neuron.titan_id_2\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5831__A1 ci_adder.uut_simple_neuron.x3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9082__CLK net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4570__A1 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7639__A2 _3621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8687__I1 ci_adder.output_memory\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4625__A2 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6910_ _3010_ _3011_ _3014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7890_ _3826_ _3830_ _3831_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_27_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6841_ _2889_ _2895_ _2950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6772_ _2806_ _2822_ _2882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8511_ ci_adder.uut_simple_neuron.x0\[11\] ci_adder.input_memory\[1\]\[11\] ci_adder.uut_simple_neuron.x2\[11\]
+ ci_adder.uut_simple_neuron.x3\[11\] _4206_ _4207_ _4219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_5723_ _1851_ _1852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5654_ _1764_ _1781_ _1784_ _1785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_45_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8442_ _4160_ _0700_ _3596_ _4161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_115_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4605_ _0740_ _0768_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8373_ ci_adder.input_memory\[1\]\[4\] _4118_ _4124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6550__A2 ci_adder.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5585_ _1699_ _1705_ _1718_ _1719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4561__A1 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7324_ _3358_ _3359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_96_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4536_ ci_adder.instruction_i\[0\] _0705_ _0687_ _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4467_ internal_ih.byte1\[2\] _0659_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7255_ _3301_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6206_ _2216_ _2215_ _2268_ _2325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_110_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7186_ ci_adder.uut_simple_neuron.titan_id_2\[20\] ci_adder.uut_simple_neuron.titan_id_5\[20\]
+ _3243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4398_ _0602_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6137_ _1958_ _2256_ _2257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_5_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ _1880_ _1997_ _2189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_84_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5019_ _1153_ _1169_ _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_68_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8709_ _0264_ net74 ci_adder.uut_simple_neuron.x3\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_36_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4552__A1 _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8294__A2 _4071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8942__CLK net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5280__I _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_17_Left_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8032__S _3908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8109__I0 internal_ih.spi_rx_byte_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _1510_ _1511_ _1512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_10_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8285__A2 _4071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7040_ ci_adder.uut_simple_neuron.titan_id_4\[28\] ci_adder.uut_simple_neuron.titan_id_3\[28\]
+ _3122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_26_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8991_ _0474_ net18 ci_adder.uut_simple_neuron.x0\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_7942_ _3703_ ci_adder.uut_simple_neuron.x2\[17\] _3855_ _3862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9249__D _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7873_ spi_interface_cvonk.SCLK_r\[2\] _3771_ _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4534__I _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout47_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6220__A1 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6824_ _2918_ _2933_ _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8815__CLK net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_35_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6755_ _2792_ _2865_ _2866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5706_ _1690_ _1809_ _1835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6686_ _2795_ _2796_ _2797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8425_ _4150_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5637_ _1766_ _1757_ _1767_ _1768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8965__CLK net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5568_ _1700_ _1702_ _1703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_8356_ spi_interface_cvonk.state\[1\] _4113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7307_ ci_adder.uut_simple_neuron.titan_id_1\[10\] ci_adder.uut_simple_neuron.titan_id_0\[10\]
+ _3344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8287_ _3625_ _4071_ _4075_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4519_ _0684_ _0688_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_41_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5499_ _1590_ _1638_ _1587_ _1639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7238_ _3264_ _3265_ _3282_ _3287_ _3288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_7169_ ci_adder.uut_simple_neuron.titan_id_2\[17\] ci_adder.uut_simple_neuron.titan_id_5\[17\]
+ ci_adder.uut_simple_neuron.titan_id_2\[16\] ci_adder.uut_simple_neuron.titan_id_5\[16\]
+ _3229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7787__A1 _3629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_53_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7539__A1 _3524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4773__A1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4380__S _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8511__I0 ci_adder.uut_simple_neuron.x0\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8027__S _3897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5253__A2 ci_adder.uut_simple_neuron.x2\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8838__CLK net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4870_ _0999_ _1024_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5005__A2 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6540_ _2592_ _2589_ _2609_ _2653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_15_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8988__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6471_ _2531_ _2568_ _2585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5422_ _1534_ _1563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8210_ ci_adder.stream_o\[31\] _3959_ _4034_ _4035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9190_ ci_adder.uut_simple_neuron.titan_id_0\[0\] net49 ci_adder.uut_simple_neuron.titan_id_2\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5353_ _1437_ _1495_ _1496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8496__I _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8141_ ci_adder.stream_o\[24\] _3959_ _3972_ _3973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5284_ _1084_ _1412_ _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8072_ _3929_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7023_ ci_adder.uut_simple_neuron.titan_id_4\[24\] ci_adder.uut_simple_neuron.titan_id_3\[24\]
+ ci_adder.uut_simple_neuron.titan_id_4\[23\] ci_adder.uut_simple_neuron.titan_id_3\[23\]
+ _3108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_65_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8974_ _0457_ net55 ci_adder.uut_simple_neuron.x0\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8164__C _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7776__S _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7925_ _3661_ ci_adder.uut_simple_neuron.x2\[9\] _3846_ _3853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7856_ internal_ih.spi_rx_byte_i\[7\] _3786_ _3784_ _3801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_38_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6807_ _2905_ _2916_ _2917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6744__A2 _2854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4999_ _0808_ _1083_ _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7787_ _3629_ _3743_ _3744_ _3745_ _3746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_6738_ _1792_ _2774_ _2849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6669_ _2723_ _2780_ _2781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__9143__CLK net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8408_ _3723_ ci_adder.input_memory\[1\]\[21\] _4139_ _4142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8339_ _4102_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_113_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9293__CLK net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7686__S _3632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4443__B1 _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout91 net92 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout80 net92 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_71_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5971_ _1919_ _2052_ _2093_ _2094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_99_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9016__CLK net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4985__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4922_ _1040_ _1073_ _1074_ _1075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7710_ _3681_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8690_ _4344_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7641_ _3455_ _3623_ _3614_ _3624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4853_ _0909_ _1007_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7923__A1 ci_adder.uut_simple_neuron.x2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9166__CLK net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4784_ _0939_ _0940_ _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4737__A1 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7572_ ci_adder.uut_simple_neuron.x0\[23\] ci_adder.uut_simple_neuron.x0\[24\] _3564_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6523_ _2632_ _2636_ _2637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_28_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9311_ _0572_ net47 ci_adder.stream_o\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9242_ _0106_ net79 ci_adder.uut_simple_neuron.titan_id_5\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6454_ _2528_ _2531_ _2568_ _2569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_113_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5405_ _1544_ _1546_ _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6385_ _2449_ _2451_ _2500_ _2501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_9173_ _0206_ net90 ci_adder.uut_simple_neuron.titan_id_3\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5336_ _1220_ _1478_ _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8124_ _3956_ _3877_ internal_ih.instruction_received _3957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5267_ _1311_ _1410_ _1411_ _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8055_ internal_ih.byte4\[7\] internal_ih.byte3\[7\] _3919_ _3921_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7006_ ci_adder.uut_simple_neuron.titan_id_4\[21\] ci_adder.uut_simple_neuron.titan_id_3\[21\]
+ _3094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6662__A1 _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5198_ _1110_ _1119_ _1343_ _1344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8957_ _0030_ net7 ci_adder.instruction_i\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7908_ _0715_ _3842_ _3844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8888_ _0435_ net32 ci_adder.output_memory\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7839_ internal_ih.spi_rx_byte_i\[2\] _3787_ _3790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7142__A2 ci_adder.uut_simple_neuron.titan_id_5\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7850__B1 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4967__A1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9189__CLK net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4719__A1 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8040__S _3908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6170_ _2244_ _2259_ _2289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5121_ _1233_ _1221_ _1268_ _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6644__A1 _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5052_ _0993_ _1133_ _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7841__B1 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8811_ _0358_ net18 internal_ih.byte3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4958__A1 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8742_ _0289_ net44 internal_ih.spi_rx_byte_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_9_Left_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5954_ _1734_ _2040_ _2077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5885_ _1945_ _1970_ _2009_ _2010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4905_ _1043_ _1058_ _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8673_ ci_adder.stream_o\[21\] ci_adder.output_memory\[21\] _4334_ _4336_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4836_ _0991_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7624_ ci_adder.normalised_stream_write_address\[1\] _0697_ _3602_ _3609_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7555_ _3540_ _3542_ _3548_ _3549_ _3550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_8_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6506_ _2047_ _2620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4767_ _0893_ _0913_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4698_ _0848_ _0857_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7486_ _3492_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6437_ _2195_ _2300_ _2552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5135__A1 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9225_ _0118_ net63 ci_adder.uut_simple_neuron.titan_id_5\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9156_ _0248_ net77 ci_adder.uut_simple_neuron.titan_id_4\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6368_ _2100_ _2249_ _2484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_101_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5319_ _1460_ _1462_ _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8107_ internal_ih.spi_rx_byte_i\[0\] _3947_ _3948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6299_ _2362_ _2369_ _2416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8475__I2 ci_adder.uut_simple_neuron.x2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9087_ _0540_ net54 ci_adder.output_val_internal\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8180__S0 _3964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8038_ internal_ih.byte3\[7\] internal_ih.byte2\[7\] _3908_ _3912_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4949__A1 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5548__I ci_adder.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7964__S _3840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7115__A2 ci_adder.uut_simple_neuron.titan_id_5\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_72_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5429__A2 _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8171__S0 _3964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4652__A3 ci_adder.uut_simple_neuron.x2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5670_ _1774_ _1776_ _1800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7729__I1 _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4621_ _0740_ _0768_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4552_ _0709_ ci_adder.uut_simple_neuron.x2\[2\] _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7340_ ci_adder.uut_simple_neuron.titan_id_1\[16\] ci_adder.uut_simple_neuron.titan_id_0\[16\]
+ _3372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7106__A2 ci_adder.uut_simple_neuron.titan_id_5\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7271_ ci_adder.uut_simple_neuron.titan_id_1\[5\] ci_adder.uut_simple_neuron.titan_id_0\[5\]
+ _3313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4483_ internal_ih.byte2\[2\] _0659_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5668__A2 _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ _2290_ _2311_ _2340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9010_ _0493_ net60 ci_adder.input_memory\[1\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6153_ _2218_ _2220_ _2272_ _2273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8162__S0 _3964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout77_I net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6084_ _2197_ _2204_ _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5104_ _1119_ _1219_ _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5035_ ci_adder.uut_simple_neuron.x2\[18\] _1184_ _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8465__S1 _4167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7968__I1 ci_adder.uut_simple_neuron.x2\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6986_ _3077_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5937_ _2038_ _2060_ _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8725_ _0280_ net25 ci_adder.uut_simple_neuron.x3\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_91_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8656_ ci_adder.stream_o\[13\] ci_adder.output_memory\[13\] _4323_ _4327_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5868_ _1963_ _1966_ _1992_ _1993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_106_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7607_ ci_adder.uut_simple_neuron.x0\[30\] ci_adder.uut_simple_neuron.x0\[31\] _3593_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_105_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5799_ _1913_ _1925_ _1926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_90_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4819_ _0973_ _0974_ _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8587_ ci_adder.uut_simple_neuron.x0\[25\] ci_adder.input_memory\[1\]\[25\] ci_adder.uut_simple_neuron.x2\[25\]
+ ci_adder.uut_simple_neuron.x3\[25\] _4252_ _4253_ _4281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_7538_ _3534_ _3535_ _3536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7469_ _3476_ _3477_ _3478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_31_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9208_ _0073_ net74 ci_adder.uut_simple_neuron.titan_id_2\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9139_ _0231_ net89 ci_adder.uut_simple_neuron.titan_id_4\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8153__S0 _3964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6608__A1 _2690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8721__CLK net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4447__I _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5831__A2 ci_adder.uut_simple_neuron.x3\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4383__S _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8871__CLK net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4570__A2 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6840_ _2940_ _2947_ _2948_ _2949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_85_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6771_ _2830_ _2840_ _2880_ _2881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5722_ _1849_ _1850_ _1851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_91_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8510_ ci_adder.output_memory\[11\] _4212_ _4218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_99_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8524__A1 _4211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5653_ _1723_ _1782_ _1783_ _1784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_5_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8441_ ci_adder.instruction_i\[0\] _0705_ _4160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7617__B _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5584_ _1686_ _1687_ _1706_ _1718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4604_ _0750_ _0751_ _0767_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8372_ _4123_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7323_ ci_adder.uut_simple_neuron.titan_id_1\[13\] ci_adder.uut_simple_neuron.titan_id_0\[13\]
+ _3358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4535_ ci_adder.instruction_i\[1\] _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6838__A1 _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4466_ _0597_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7254_ ci_adder.uut_simple_neuron.titan_id_2\[31\] ci_adder.uut_simple_neuron.titan_id_5\[31\]
+ _3300_ _3301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_6205_ _2165_ _2117_ _2164_ _2160_ _2219_ _2324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_68_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7185_ _3242_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4397_ _0622_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6136_ _1960_ _2097_ _2256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_5_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6067_ _2137_ _2186_ _2187_ _2188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8894__CLK net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5018_ _1155_ _1168_ _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_68_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8602__I2 _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5577__A1 _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6969_ ci_adder.uut_simple_neuron.titan_id_4\[15\] ci_adder.uut_simple_neuron.titan_id_3\[15\]
+ _3063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8708_ _0263_ net81 ci_adder.uut_simple_neuron.x3\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__8515__A1 ci_adder.output_memory\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8639_ ci_adder.stream_o\[5\] ci_adder.output_memory\[5\] _4312_ _4318_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_106_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5568__A1 _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7801__I0 _3757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8313__S _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8109__I1 internal_ih.current_instruction\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8767__CLK net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input1_I spi_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8990_ _0473_ net25 ci_adder.uut_simple_neuron.x0\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_7941_ _3861_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7872_ _3812_ _3815_ _3816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_38_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5559__A1 _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6823_ _2921_ _2932_ _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6754_ _2794_ _2864_ _2865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6685_ _2767_ _2778_ _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5705_ _1795_ _1832_ _1833_ _1834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_98_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout6_I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5636_ _1750_ _1756_ _1767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8424_ _3762_ ci_adder.input_memory\[1\]\[29\] _4139_ _4150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7720__A2 _3659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5567_ _1679_ _1701_ _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_4
X_8355_ _3786_ _3780_ _4112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ _1544_ _1546_ _1586_ _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7306_ _3343_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4518_ ci_adder.instruction_i\[0\] ci_adder.instruction_i\[1\] _0687_ _0688_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8286_ ci_adder.uut_simple_neuron.x0\[2\] _4072_ _4075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7237_ ci_adder.uut_simple_neuron.titan_id_2\[27\] ci_adder.uut_simple_neuron.titan_id_5\[27\]
+ _3281_ _3284_ _3286_ _3287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4449_ _0650_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7168_ _3221_ _3226_ _3228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6119_ _1919_ _2049_ _2239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7099_ _3169_ _3170_ _3171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_107_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9072__CLK net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6278__A2 _2349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5789__A1 ci_adder.uut_simple_neuron.x3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7778__A2 _3659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5253__A3 ci_adder.uut_simple_neuron.x2\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_15_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6470_ _2531_ _2568_ _2584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5713__A1 ci_adder.uut_simple_neuron.x3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5421_ _1528_ _1535_ _1561_ _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5352_ _1494_ _1495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8140_ _3960_ _3969_ _3971_ _3815_ _3972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_23_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8071_ internal_ih.byte5\[7\] internal_ih.byte4\[7\] _3919_ _3929_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7022_ _3100_ _3105_ _3107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5283_ _1392_ _1425_ _1426_ _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4545__I _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8973_ _0456_ net60 ci_adder.uut_simple_neuron.x0\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_78_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7924_ _3654_ _3842_ _3852_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7855_ _3770_ _3799_ _3800_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6806_ _2908_ _2915_ _2916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4998_ _1116_ _1147_ _1148_ _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7786_ ci_adder.value_i\[26\] _3608_ _3745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6737_ _1801_ _1810_ _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8577__S0 _4252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6668_ _2766_ _2779_ _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6599_ _2706_ _2711_ _2712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5619_ ci_adder.uut_simple_neuron.x3\[5\] ci_adder.uut_simple_neuron.x3\[6\] _1751_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_61_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8407_ _4141_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8338_ _3751_ ci_adder.uut_simple_neuron.x0\[27\] _4091_ _4102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8269_ ci_adder.uut_simple_neuron.titan_id_6\[28\] _4065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_113_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4691__A1 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4443__B2 internal_ih.byte2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout92 net4 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout81 net84 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout70 net92 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_12_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7448__A1 ci_adder.uut_simple_neuron.x0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6120__A1 _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8805__CLK net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8038__S _3908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8955__CLK net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5970_ _2049_ _2051_ _2093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_87_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4921_ _1044_ _1061_ _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6187__A1 _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4852_ _0894_ _0975_ _1006_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8420__I0 _3751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7640_ ci_adder.uut_simple_neuron.x0\[0\] ci_adder.uut_simple_neuron.x0\[1\] ci_adder.uut_simple_neuron.x0\[2\]
+ _3623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__7923__A2 _3846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4783_ _0928_ _0909_ _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_74_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_72_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7571_ _3561_ _3562_ _3563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6522_ _2634_ _2635_ _2636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9310_ _0571_ net47 ci_adder.stream_o\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6453_ _2557_ _2567_ _2568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9241_ _0105_ net75 ci_adder.uut_simple_neuron.titan_id_5\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5404_ _0996_ _1499_ _1545_ _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9172_ _0205_ net88 ci_adder.uut_simple_neuron.titan_id_3\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6384_ _2458_ _2460_ _2499_ _2500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8123_ net12 _3956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_100_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5335_ ci_adder.uut_simple_neuron.x2\[23\] _1267_ _1398_ _1478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5266_ _1310_ _1357_ _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8054_ _3920_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7005_ _3093_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5197_ _1340_ _1341_ _1342_ _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_97_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8956_ _0029_ net7 ci_adder.instruction_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7907_ _3616_ _3841_ _3843_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4425__B2 internal_ih.byte1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6178__A1 _2249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8887_ _0434_ net35 ci_adder.output_memory\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9110__CLK net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7838_ internal_ih.spi_tx_byte_o\[1\] _3779_ _3784_ internal_ih.spi_rx_byte_i\[1\]
+ _3789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_93_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5925__A1 ci_adder.uut_simple_neuron.x3\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7769_ ci_adder.uut_simple_neuron.x0\[23\] _3726_ _3731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7678__A1 ci_adder.uut_simple_neuron.x3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9260__CLK net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8828__CLK net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6653__A2 _2764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4386__S _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4664__A1 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_126_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4416__B2 internal_ih.byte1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4967__A2 _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7669__A1 _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_77_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6341__A1 _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5120_ _1233_ ci_adder.uut_simple_neuron.x2\[22\] _1268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5051_ _1141_ _1199_ _1201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4407__A1 internal_ih.byte4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8810_ _0357_ net18 internal_ih.byte3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9133__CLK net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8741_ _0288_ net44 internal_ih.spi_rx_byte_i\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4407__B2 internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5953_ _2035_ _2061_ _2075_ _2076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_88_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4958__A2 _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5080__A1 _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5884_ _1947_ _1969_ _2009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_80_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4904_ _1056_ _1057_ _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_8_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8672_ _4335_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5907__A1 _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4835_ _0989_ _0990_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_63_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7623_ _3604_ _3608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_fanout22_I net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ _0896_ _0912_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7554_ ci_adder.uut_simple_neuron.x0\[19\] ci_adder.uut_simple_neuron.x0\[21\] _3539_
+ _3549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6505_ _2617_ _2618_ _2619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4697_ _0849_ _0856_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7485_ _3488_ _3491_ _3492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6436_ _2535_ _2548_ _2550_ _2551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_31_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9224_ _0107_ net50 ci_adder.uut_simple_neuron.titan_id_5\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9155_ _0247_ net76 ci_adder.uut_simple_neuron.titan_id_4\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6367_ _2466_ _2482_ _2483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5318_ _0996_ _1416_ _1461_ _1462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4894__A1 _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8106_ _3816_ _3818_ _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_110_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6298_ _2371_ _2415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8475__I3 ci_adder.uut_simple_neuron.x3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9086_ _0539_ net34 ci_adder.output_val_internal\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5249_ _1344_ _1360_ _1393_ _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8037_ _3911_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8406__S _4139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_119_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8939_ _0003_ net8 ci_adder.address_i\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4885__A1 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7823__A1 _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8379__A2 _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5062__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4620_ _0742_ _0773_ _0775_ _0765_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__8551__A2 _4212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4551_ _0710_ _0718_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8303__A2 _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6314__A1 _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7270_ _3312_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4482_ _0667_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6221_ _2290_ _2311_ _2339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6152_ _2162_ _2160_ _2215_ _2272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_0_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5103_ _1151_ _1219_ _1250_ _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6083_ _2051_ _2203_ _2204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4628__A1 _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5034_ ci_adder.uut_simple_neuron.x2\[19\] ci_adder.uut_simple_neuron.x2\[20\] _1184_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_79_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6985_ _3075_ _3076_ _3077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5936_ _2042_ _2059_ _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4800__A1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8724_ _0279_ net25 ci_adder.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_8655_ _4326_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ _1956_ _1962_ _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8542__A2 _4243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7606_ _3590_ _3591_ _3592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6553__A1 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5798_ _1922_ _1924_ _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4818_ ci_adder.uut_simple_neuron.x2\[12\] ci_adder.uut_simple_neuron.x2\[13\] ci_adder.uut_simple_neuron.x2\[14\]
+ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_8_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8586_ ci_adder.output_memory\[25\] _4258_ _4280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4749_ ci_adder.uut_simple_neuron.x2\[9\] _0905_ _0906_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7537_ ci_adder.uut_simple_neuron.x0\[18\] ci_adder.uut_simple_neuron.x0\[19\] _3535_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6305__A1 _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7468_ _3469_ _3470_ _3477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6419_ _2470_ _2478_ _2534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_9207_ _0072_ net84 ci_adder.uut_simple_neuron.titan_id_2\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9179__CLK net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7399_ _3415_ _3418_ _3419_ _3420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9138_ _0230_ net87 ci_adder.uut_simple_neuron.titan_id_4\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9069_ _0522_ net61 ci_adder.output_val_internal\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5292__A1 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5044__A1 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8533__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8297__A1 _3470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4858__A1 _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8696__CLK net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8046__S _3908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5035__A1 ci_adder.uut_simple_neuron.x2\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6770_ _2804_ _2828_ _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6783__A1 ci_adder.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5721_ _1702_ _1752_ _1850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_85_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6535__A1 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ _1748_ _1758_ _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8440_ _3974_ _4158_ _4159_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5583_ _1678_ _1716_ _1717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4603_ ci_adder.uut_simple_neuron.x2\[2\] ci_adder.uut_simple_neuron.x2\[5\] _0767_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_60_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8371_ _3631_ ci_adder.input_memory\[1\]\[3\] _4122_ _4123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7322_ ci_adder.uut_simple_neuron.titan_id_1\[12\] ci_adder.uut_simple_neuron.titan_id_0\[12\]
+ _3354_ _3355_ _3357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_53_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9321__CLK net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4534_ _0703_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XTAP_TAPCELL_ROW_96_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4465_ _0658_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7253_ _3296_ _3297_ _3299_ _3300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6204_ _2322_ _2271_ _2323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7184_ _3240_ _3241_ _3242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4396_ internal_ih.byte4\[1\] _0603_ _0620_ internal_ih.byte0\[1\] _0622_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6135_ _2247_ _2254_ _2255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6066_ _2139_ _2152_ _2187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5017_ _1157_ _1167_ _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8063__I1 internal_ih.byte4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8602__I3 ci_adder.uut_simple_neuron.x3\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6968_ _3062_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8707_ _0262_ net81 ci_adder.uut_simple_neuron.x3\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_52_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5919_ _1880_ _2000_ _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6899_ ci_adder.uut_simple_neuron.titan_id_4\[3\] ci_adder.uut_simple_neuron.titan_id_3\[3\]
+ _3005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_64_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8515__A2 _4212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8638_ _4317_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8569_ ci_adder.output_val_internal\[21\] _4249_ _4267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7254__A2 ci_adder.uut_simple_neuron.titan_id_5\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7801__I1 ci_adder.uut_simple_neuron.x3\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5568__A2 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7718__B ci_adder.uut_simple_neuron.x0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7940_ _3697_ ci_adder.uut_simple_neuron.x2\[16\] _3855_ _3861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7871_ _3807_ _3808_ _3814_ _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_TAPCELL_ROW_38_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6822_ _2924_ _2931_ _2932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5559__A2 _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6753_ _2859_ _2863_ _2864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6684_ _2768_ _2769_ _2777_ _2795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5704_ _1799_ _1812_ _1833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5635_ _1750_ _1756_ _1766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8423_ _4149_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8711__CLK net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5566_ ci_adder.uut_simple_neuron.x3\[3\] ci_adder.uut_simple_neuron.x3\[4\] _1701_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8354_ spi_interface_cvonk.state\[1\] spi_interface_cvonk.state\[0\] _4111_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5497_ _1596_ _1636_ _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7305_ _3341_ _3342_ _3343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4517_ ci_adder.instruction_i\[2\] _0685_ _0686_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8285_ _3621_ _4071_ _4074_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7236_ _3285_ _3286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4448_ internal_ih.byte0\[1\] _0648_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_1_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7167_ _3227_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4379_ _0610_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6118_ _2192_ _2236_ _2237_ _2238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5247__A1 _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7098_ ci_adder.uut_simple_neuron.titan_id_2\[6\] ci_adder.uut_simple_neuron.titan_id_5\[6\]
+ _3170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6049_ _2122_ _2155_ _2170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_107_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8036__I1 internal_ih.byte2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8587__I2 ci_adder.uut_simple_neuron.x2\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8197__B1 ci_adder.stream_o\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8414__S _4139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5970__A2 _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4389__S _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5789__A2 ci_adder.uut_simple_neuron.x3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8324__S _4091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8123__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5713__A2 ci_adder.uut_simple_neuron.x3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5420_ _1525_ _1537_ _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5351_ _1475_ _1493_ _1494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5282_ _1394_ _1414_ _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8070_ _3928_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7021_ _3106_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8972_ _0455_ net55 ci_adder.uut_simple_neuron.x0\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_7923_ ci_adder.uut_simple_neuron.x2\[8\] _3846_ _3852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout52_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7854_ internal_ih.spi_rx_byte_i\[7\] _3787_ _3800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6805_ _2914_ _2915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7785_ ci_adder.uut_simple_neuron.x0\[26\] _3562_ _3730_ _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_108_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6736_ _2845_ _2846_ _2847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_102_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4997_ _1118_ _1130_ _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8577__S1 _4253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6667_ _2767_ _2778_ _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_18_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6598_ _2517_ _2707_ _2710_ _2711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5618_ _1692_ _1733_ _1749_ _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_8406_ _3718_ ci_adder.input_memory\[1\]\[20\] _4139_ _4141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5549_ _1684_ _1676_ _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8337_ _4101_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8268_ _4064_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_113_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7219_ _3269_ _3271_ _3272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8199_ _3811_ _4024_ _4025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_100_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5640__A1 _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout71 net72 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout82 net83 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout60 net70 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_52_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7940__I0 _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7448__A2 _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4646__I _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4920_ _1044_ _1061_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4851_ _0899_ ci_adder.uut_simple_neuron.x2\[13\] ci_adder.uut_simple_neuron.x2\[14\]
+ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_51_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4782_ _0904_ _0937_ _0938_ _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_55_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7570_ ci_adder.uut_simple_neuron.x0\[24\] ci_adder.uut_simple_neuron.x0\[25\] _3562_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ _1750_ _1757_ _2635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6452_ _2560_ _2566_ _2567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9240_ _0104_ net74 ci_adder.uut_simple_neuron.titan_id_5\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5403_ _1467_ _1498_ _1545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_9171_ _0204_ net88 ci_adder.uut_simple_neuron.titan_id_3\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9062__CLK net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6101__I _2221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6383_ _2462_ _2488_ _2498_ _2499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_101_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8122_ _3955_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5334_ _0717_ _1449_ _1448_ _1476_ _1402_ _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_5265_ _1310_ _1357_ _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8053_ internal_ih.byte4\[6\] internal_ih.byte3\[6\] _3919_ _3920_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7641__B _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7004_ _3091_ _3092_ _3093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5196_ _1310_ _1313_ _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5870__A1 _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4673__A2 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7998__I0 internal_ih.byte1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5622__A1 ci_adder.uut_simple_neuron.x3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4425__A2 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8955_ _0028_ net11 ci_adder.instruction_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7906_ _0710_ _3842_ _3843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8886_ _0433_ net34 ci_adder.output_memory\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7837_ _3770_ _3785_ _3788_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8191__C _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7768_ ci_adder.uut_simple_neuron.x0\[23\] _3726_ _3730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6719_ _2829_ _2830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7699_ _3672_ ci_adder.uut_simple_neuron.x3\[11\] _3632_ _3673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7678__A2 _3617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_115_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4466__I _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8650__I1 ci_adder.output_memory\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4416__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7669__A2 _3470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7913__I0 _3631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6341__A2 _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8618__A1 _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8922__CLK net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5050_ _1142_ _1199_ _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8641__I1 ci_adder.output_memory\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5952_ _2038_ _2060_ _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5604__A1 _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8740_ _0287_ net42 internal_ih.spi_rx_byte_i\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4407__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4903_ _1011_ ci_adder.uut_simple_neuron.x2\[16\] _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5883_ _1985_ _1987_ _2007_ _2008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_118_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8671_ ci_adder.stream_o\[20\] ci_adder.output_memory\[20\] _4334_ _4335_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4834_ _0950_ _0948_ _0988_ _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_75_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7622_ _3603_ _3606_ _3607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_117_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4765_ _0804_ _0915_ _0921_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7553_ _3539_ ci_adder.uut_simple_neuron.x0\[21\] _3548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6504_ _1734_ _2564_ _2618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4696_ _0713_ _0850_ _0855_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_70_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7484_ _3489_ _3490_ _3491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_9223_ _0096_ net50 ci_adder.uut_simple_neuron.titan_id_5\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6435_ _2199_ _2549_ _2550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9154_ _0246_ net76 ci_adder.uut_simple_neuron.titan_id_4\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6366_ _2479_ _2481_ _2482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5317_ _1389_ _1415_ _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8105_ _3946_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9085_ _0538_ net34 ci_adder.output_val_internal\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6297_ _2362_ _2369_ _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8036_ internal_ih.byte3\[6\] internal_ih.byte2\[6\] _3908_ _3911_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_110_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5248_ _1346_ _1359_ _1393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5179_ _1281_ _1284_ _1326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8938_ _0002_ net8 ci_adder.address_i\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8869_ _0416_ net50 ci_adder.output_memory\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_121_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8422__S _4139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6020__A1 _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4582__A1 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8945__CLK net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6676__I _2787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8320__I0 _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5834__A1 ci_adder.uut_simple_neuron.x3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8387__I0 _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8332__S _4091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4573__A1 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4550_ _0717_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_107_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ internal_ih.byte2\[1\] _0659_ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_123_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6220_ _1695_ _2337_ _2338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6151_ _2268_ _2270_ _2271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6078__A1 _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5102_ _1084_ _1218_ _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5825__A1 _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6082_ _2199_ _2202_ _2203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5033_ _0711_ _1163_ _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6250__A1 _2364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6984_ ci_adder.uut_simple_neuron.titan_id_4\[18\] ci_adder.uut_simple_neuron.titan_id_3\[18\]
+ _3076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8818__CLK net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5935_ _2045_ _2058_ _2059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8723_ _0278_ net28 ci_adder.uut_simple_neuron.x3\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5866_ _1709_ _1990_ _1991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_76_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8654_ ci_adder.stream_o\[12\] ci_adder.output_memory\[12\] _4323_ _4326_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6002__A1 _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4817_ _0899_ ci_adder.uut_simple_neuron.x2\[13\] ci_adder.uut_simple_neuron.x2\[14\]
+ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7605_ _3585_ _3588_ _3591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5797_ _1730_ _1923_ _1924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8968__CLK net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8585_ _4257_ _4276_ _4278_ _4279_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_105_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4564__A1 _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4748_ ci_adder.uut_simple_neuron.x2\[10\] ci_adder.uut_simple_neuron.x2\[11\] _0906_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7536_ ci_adder.uut_simple_neuron.x0\[18\] ci_adder.uut_simple_neuron.x0\[19\] _3534_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4679_ _0832_ _0839_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7467_ _3459_ _3469_ _3476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6418_ _2483_ _2487_ _2532_ _2533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9206_ _0071_ net81 ci_adder.uut_simple_neuron.titan_id_2\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9137_ _0229_ net87 ci_adder.uut_simple_neuron.titan_id_4\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7398_ ci_adder.uut_simple_neuron.titan_id_1\[26\] ci_adder.uut_simple_neuron.titan_id_0\[26\]
+ _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6349_ _2420_ _2426_ _2465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6069__A1 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9068_ _0521_ net48 ci_adder.output_val_internal\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7805__A2 _3629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8019_ internal_ih.byte2\[6\] internal_ih.byte1\[6\] _3897_ _3902_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8297__A2 _4072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8541__I0 _3524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9123__CLK net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4858__A2 ci_adder.uut_simple_neuron.x2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5720_ _1700_ _1849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5651_ _1748_ _1758_ _1782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7732__A1 _3524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5582_ _1709_ _1715_ _1716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4602_ ci_adder.uut_simple_neuron.x2\[6\] _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8370_ _4116_ _4122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7321_ _3356_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4533_ ci_adder.address_i\[2\] _0702_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_96_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7252_ ci_adder.uut_simple_neuron.titan_id_2\[30\] ci_adder.uut_simple_neuron.titan_id_5\[30\]
+ _3299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_41_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6203_ _2215_ _2217_ _2322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_123_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4849__A2 _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4464_ internal_ih.byte1\[1\] _0648_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7183_ ci_adder.uut_simple_neuron.titan_id_2\[20\] ci_adder.uut_simple_neuron.titan_id_5\[20\]
+ _3241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4395_ _0621_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6134_ _2100_ _2253_ _2254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_0_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6065_ _2139_ _2152_ _2186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_5_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5016_ _1158_ _1166_ _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6967_ ci_adder.uut_simple_neuron.titan_id_4\[15\] ci_adder.uut_simple_neuron.titan_id_3\[15\]
+ _3061_ _3062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5918_ _1728_ _2041_ _2042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_105_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8706_ _0261_ net81 ci_adder.uut_simple_neuron.x3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_52_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6898_ ci_adder.uut_simple_neuron.titan_id_4\[3\] ci_adder.uut_simple_neuron.titan_id_3\[3\]
+ _3004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_36_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5849_ _1971_ _1974_ _1975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8637_ ci_adder.stream_o\[4\] ci_adder.output_memory\[4\] _4312_ _4317_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9146__CLK net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4537__A1 _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8568_ _4260_ _4265_ _4266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7519_ _3508_ ci_adder.uut_simple_neuron.x0\[15\] _3520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8499_ _4165_ _4208_ _4209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6765__A2 _2854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4776__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7962__A1 _3751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7714__A1 _3619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8057__S _3919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9019__CLK net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7870_ internal_ih.instruction_received internal_ih.spi_rx_byte_i\[3\] _3813_ _3814_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6821_ _0163_ _2930_ _2931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5559__A3 _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7953__A1 _3728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6752_ _2861_ _2862_ _2863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9169__CLK net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6683_ _2793_ _2784_ _2794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5703_ _1799_ _1812_ _1832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5634_ _1677_ _1700_ _1765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_72_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8422_ _3757_ ci_adder.input_memory\[1\]\[28\] _4139_ _4149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8353_ spi_interface_cvonk.state\[0\] _4109_ _4110_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5565_ _1676_ _1691_ _1687_ _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7304_ ci_adder.uut_simple_neuron.titan_id_1\[10\] ci_adder.uut_simple_neuron.titan_id_0\[10\]
+ _3342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5496_ _0996_ _1635_ _1636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4516_ ci_adder.instruction_i\[4\] ci_adder.instruction_i\[7\] ci_adder.instruction_i\[6\]
+ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_8284_ ci_adder.uut_simple_neuron.x0\[1\] _4072_ _4074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7235_ ci_adder.uut_simple_neuron.titan_id_2\[27\] ci_adder.uut_simple_neuron.titan_id_5\[27\]
+ ci_adder.uut_simple_neuron.titan_id_2\[26\] ci_adder.uut_simple_neuron.titan_id_5\[26\]
+ _3285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4447_ _0649_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7166_ _3225_ _3226_ _3227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6117_ _2194_ _2209_ _2237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_13_Left_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4378_ internal_ih.byte7\[3\] _0603_ _0609_ net14 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6444__A1 _1715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7097_ _3165_ _3168_ _3169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6048_ _2169_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_107_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7944__A1 _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8587__I3 ci_adder.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7999_ _3891_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4758__A1 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8511__I3 ci_adder.uut_simple_neuron.x3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_69_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9311__CLK net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8340__S _4070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5350_ _1400_ _1492_ _1493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_93_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5281_ _1394_ _1414_ _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7020_ _3104_ _3105_ _3106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8971_ _0454_ net58 ci_adder.uut_simple_neuron.x0\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4437__B1 _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7922_ _3650_ _3842_ _3851_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7853_ internal_ih.spi_tx_byte_o\[6\] _3779_ _3784_ internal_ih.spi_rx_byte_i\[6\]
+ _3799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_fanout45_I net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6804_ _2911_ _2913_ _2914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4996_ _1118_ _1130_ _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7784_ _3562_ _3730_ ci_adder.uut_simple_neuron.x0\[26\] _3743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6735_ _2757_ _2763_ _2846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_102_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6666_ _2770_ _2777_ _2778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6597_ _2708_ _2579_ _2709_ _2710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5617_ _1730_ _1732_ _1749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8405_ _4140_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5548_ ci_adder.uut_simple_neuron.x3\[0\] _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_60_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8336_ _3746_ ci_adder.uut_simple_neuron.x0\[26\] _4091_ _4101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8267_ ci_adder.uut_simple_neuron.titan_id_6\[27\] _4064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5479_ _1573_ _1618_ _1619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7218_ _3264_ _3265_ _3270_ _3271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_113_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8198_ ci_adder.output_val_internal\[30\] ci_adder.output_val_internal\[22\] ci_adder.output_val_internal\[14\]
+ ci_adder.output_val_internal\[6\] _3964_ _3961_ _4024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7149_ ci_adder.uut_simple_neuron.titan_id_2\[14\] ci_adder.uut_simple_neuron.titan_id_5\[14\]
+ _3213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5640__A2 _1754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7917__A1 ci_adder.uut_simple_neuron.x2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout83 net84 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout72 net80 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_64_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout61 net69 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_12_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout50 net51 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_64_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5156__A1 _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4903__A1 _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7940__I1 ci_adder.uut_simple_neuron.x2\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7853__B1 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7908__A1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4850_ _0939_ _0967_ _1004_ _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8134__I _3964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8851__CLK net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8581__A1 ci_adder.output_memory\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6520_ _1723_ _2633_ _2634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4781_ _0936_ _0907_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_28_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6451_ _2563_ _2565_ _2566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6382_ _2491_ _2497_ _2498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5402_ _0994_ _1543_ _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9170_ _0203_ net89 ci_adder.uut_simple_neuron.titan_id_3\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5333_ _1451_ _1476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8121_ internal_ih.current_instruction\[7\] _3947_ _3955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5264_ _1397_ _1408_ _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8052_ _3818_ _3919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7844__B1 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7003_ ci_adder.uut_simple_neuron.titan_id_4\[21\] ci_adder.uut_simple_neuron.titan_id_3\[21\]
+ _3092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5195_ _1310_ _1313_ _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4673__A3 ci_adder.uut_simple_neuron.x2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7998__I1 internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8954_ _0027_ net10 ci_adder.instruction_i\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7905_ _3840_ _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8885_ _0432_ net34 ci_adder.output_memory\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7836_ internal_ih.spi_rx_byte_i\[1\] _3787_ _3788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4979_ _1118_ _1130_ _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7767_ _3617_ _3728_ _3729_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6718_ _2804_ _2828_ _2829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7127__A2 ci_adder.uut_simple_neuron.titan_id_5\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7698_ _3629_ _3669_ _3670_ _3671_ _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_117_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6649_ _2190_ _2207_ _2761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_115_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8319_ _4092_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9299_ _0560_ net49 ci_adder.stream_o\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8724__CLK net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_126_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6810__A1 _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8874__CLK net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7118__A2 ci_adder.uut_simple_neuron.titan_id_5\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5129__A1 _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7913__I1 _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8618__A2 _4305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5301__A1 ci_adder.uut_simple_neuron.x2\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8065__S _3919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5951_ _2023_ _2064_ _2074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_88_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ _1011_ _1055_ _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8670_ _3601_ _4334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5882_ _1991_ _1993_ _2006_ _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_75_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4833_ _0950_ _0948_ _0988_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7621_ _3604_ _3605_ _3606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4764_ _0879_ _0914_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7552_ ci_adder.uut_simple_neuron.x0\[21\] ci_adder.uut_simple_neuron.x0\[22\] _3547_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6503_ _2040_ _2056_ _2617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7483_ _3470_ ci_adder.uut_simple_neuron.x0\[9\] _3479_ _3490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_15_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6434_ _2202_ _2364_ _2549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4695_ _0851_ _0854_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9222_ ci_adder.uut_simple_neuron.titan_id_3\[0\] net49 ci_adder.uut_simple_neuron.titan_id_5\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9153_ _0245_ net76 ci_adder.uut_simple_neuron.titan_id_4\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6365_ _2143_ _2480_ _2481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8747__CLK net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8609__A2 _4161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6296_ _2357_ _2411_ _2412_ _2413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5316_ _0993_ _1459_ _1460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8104_ internal_ih.byte7\[7\] internal_ih.byte6\[7\] _3825_ _3946_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9084_ _0537_ net54 ci_adder.output_val_internal\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5247_ _1151_ _1390_ _1391_ _1392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8035_ _3910_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_110_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8897__CLK net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5178_ _0996_ _1293_ _1324_ _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_79_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8937_ _0024_ net9 ci_adder.address_i\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8868_ _0415_ net63 ci_adder.output_memory\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5359__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7819_ spi_interface_cvonk.SCLK_r\[2\] _3771_ _3772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8799_ _0346_ net22 internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_121_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6020__A2 _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8502__I _4161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5531__A1 ci_adder.uut_simple_neuron.x2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5598__A1 ci_adder.uut_simple_neuron.x3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9052__CLK net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4573__A2 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4480_ _0666_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6150_ _2216_ _2215_ _2269_ _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5101_ _1217_ _1238_ _1239_ _1156_ _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_0_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6081_ _2098_ _2201_ _2202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5825__A2 _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5032_ _0718_ _1181_ _1165_ _1159_ _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5589__A1 _1721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6983_ _3073_ _3074_ _3075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_69_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5934_ _2054_ _2057_ _2058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8722_ _0277_ net72 ci_adder.uut_simple_neuron.x3\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5865_ _1715_ _1989_ _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8653_ _4325_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4816_ _0970_ _0971_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_76_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7604_ ci_adder.uut_simple_neuron.x0\[29\] ci_adder.uut_simple_neuron.x0\[30\] _3590_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5796_ _1732_ _1803_ _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8584_ ci_adder.output_val_internal\[24\] _4249_ _4279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4564__A2 ci_adder.uut_simple_neuron.x2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4747_ ci_adder.uut_simple_neuron.x2\[10\] ci_adder.uut_simple_neuron.x2\[11\] _0905_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7535_ _3532_ _3533_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4678_ _0833_ _0838_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7466_ _3465_ _3466_ _3474_ _3464_ _3475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_31_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6417_ _2466_ _2482_ _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9205_ _0070_ net82 ci_adder.uut_simple_neuron.titan_id_2\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7397_ ci_adder.uut_simple_neuron.titan_id_1\[26\] ci_adder.uut_simple_neuron.titan_id_0\[26\]
+ _3418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6348_ _2428_ _2464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_101_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9136_ _0228_ net91 ci_adder.uut_simple_neuron.titan_id_4\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8138__S0 _3964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6279_ _2344_ _2350_ _2396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9067_ _0520_ net61 ci_adder.output_val_internal\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8018_ _3901_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8912__CLK net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5752__A1 ci_adder.uut_simple_neuron.x3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4858__A3 ci_adder.uut_simple_neuron.x2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8206__B1 ci_adder.stream_o\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6232__A2 _2349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8509__A1 _4211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5650_ _1765_ _1780_ _1781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4670__I _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4601_ _0763_ _0764_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_26_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5581_ _1681_ _1714_ _1715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5743__A1 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7320_ _3354_ _3355_ _3356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4532_ _0696_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4463_ _0657_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7251_ _3298_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6202_ _2318_ _2320_ _2321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_123_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7182_ _3238_ _3239_ _3240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4394_ internal_ih.byte4\[0\] _0603_ _0620_ internal_ih.byte0\[0\] _0621_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__9098__CLK net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6133_ _2249_ _2252_ _2253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6064_ _2126_ _2184_ _2185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout75_I net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7799__A2 _3659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_77_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5015_ _1159_ _1165_ _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8048__I0 internal_ih.byte4\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8317__I _4070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6966_ _3057_ _3058_ _3060_ _3061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5917_ _1734_ _2040_ _2041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8705_ _0260_ net82 ci_adder.uut_simple_neuron.x3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_52_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5982__A1 _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6897_ _3003_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8052__I _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _1972_ _1973_ _1974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8636_ _4316_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5779_ _1872_ _1889_ _1905_ _1906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_86_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8567_ ci_adder.uut_simple_neuron.x0\[21\] ci_adder.input_memory\[1\]\[21\] _1233_
+ _2365_ _4252_ _4253_ _4265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_32_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7518_ _3510_ _3511_ _3518_ _3509_ _3519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_44_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8498_ ci_adder.uut_simple_neuron.x0\[9\] ci_adder.input_memory\[1\]\[9\] ci_adder.uut_simple_neuron.x2\[9\]
+ ci_adder.uut_simple_neuron.x3\[9\] _4206_ _4207_ _4208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_101_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7449_ _3453_ _3457_ _3461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9119_ _0184_ net27 ci_adder.uut_simple_neuron.titan_id_0\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8428__S _4116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_95_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8531__S0 _4206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4473__A1 internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7962__A2 _3846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A1 ci_adder.uut_simple_neuron.x3\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7478__A1 _3479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9240__CLK net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8808__CLK net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8338__S _4091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8958__CLK net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6820_ _2927_ _2929_ _2930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7953__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6751_ _2720_ _2781_ _2862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6682_ _2720_ _2781_ _2793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5702_ _1828_ _1816_ _1830_ _1831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5633_ _1763_ _1759_ _1764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5716__A1 ci_adder.uut_simple_neuron.x3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8421_ _4148_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5564_ _1690_ _1697_ _1698_ _1699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8352_ _3786_ _3780_ spi_interface_cvonk.state\[0\] _4110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7303_ _3337_ _3339_ _3340_ _3341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_5_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4515_ ci_adder.instruction_i\[3\] ci_adder.instruction_i\[5\] _0685_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5495_ _1599_ _1634_ _1635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8283_ _3616_ _4071_ _4073_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7234_ _3270_ _3283_ _3268_ _3284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4446_ internal_ih.byte0\[0\] _0648_ _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7165_ ci_adder.uut_simple_neuron.titan_id_2\[17\] ci_adder.uut_simple_neuron.titan_id_5\[17\]
+ _3226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4377_ internal_ih.byte4\[3\] internal_ih.byte3\[3\] _0599_ _0609_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6116_ _2194_ _2209_ _2236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4575__I _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7096_ _3166_ _3167_ _3168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6047_ _2164_ _2168_ _2169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_107_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7944__A2 _3846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9113__CLK net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7998_ internal_ih.byte1\[4\] internal_ih.byte0\[4\] _3886_ _3891_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6949_ ci_adder.uut_simple_neuron.titan_id_4\[11\] ci_adder.uut_simple_neuron.titan_id_3\[11\]
+ _3047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8619_ ci_adder.output_val_internal\[31\] _4161_ _4307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_118_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6380__A1 _1715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8121__A2 _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6132__A1 ci_adder.uut_simple_neuron.x3\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4446__A1 internal_ih.byte0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8188__A2 ci_adder.stream_o\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7745__B _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8112__A2 _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5280_ _1424_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_93_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8780__CLK net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8970_ _0453_ net58 ci_adder.uut_simple_neuron.x0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__9136__CLK net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7921_ _0787_ _3846_ _3851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4437__B2 internal_ih.byte2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8179__A2 ci_adder.stream_o\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7852_ _3770_ _3797_ _3798_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6803_ _1882_ _2912_ _2913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4995_ _0993_ _1133_ _1145_ _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7783_ _3742_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout38_I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9286__CLK net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6734_ _2760_ _2762_ _2845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_102_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6665_ _1675_ _2776_ _2777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7154__A3 _3216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8404_ _3713_ ci_adder.input_memory\[1\]\[19\] _4139_ _4140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6596_ _2643_ _2709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5616_ _1725_ _1746_ _1747_ _1748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_104_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5547_ _1683_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8335_ _4100_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5478_ _1614_ _1617_ _1618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8266_ _4063_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7217_ ci_adder.uut_simple_neuron.titan_id_2\[24\] ci_adder.uut_simple_neuron.titan_id_5\[24\]
+ _3270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4429_ internal_ih.byte6\[0\] _0635_ _0632_ internal_ih.byte2\[0\] _0640_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7862__A1 internal_ih.spi_rx_byte_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4676__A1 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8197_ _3963_ ci_adder.stream_o\[6\] ci_adder.stream_o\[22\] _3965_ _4022_ _4023_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_7148_ _3208_ _3210_ _3211_ _3212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7079_ _3153_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7090__A2 ci_adder.uut_simple_neuron.titan_id_5\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8414__I0 _3736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8505__I _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7917__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout40 net92 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4600__A1 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout73 net75 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout62 net69 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_12_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout51 net52 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout84 net90 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4903__A2 ci_adder.uut_simple_neuron.x2\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9009__CLK net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9159__CLK net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7908__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5919__A1 _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4780_ _0936_ _0907_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_28_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6450_ _1734_ _2564_ _2565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_125_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6381_ _2494_ _2496_ _2497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5401_ _1516_ _1542_ _1543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ _1400_ _1453_ _1474_ _1475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_51_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8120_ _3954_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4658__A1 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5263_ _1400_ _1407_ _1408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7844__B2 internal_ih.spi_rx_byte_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8051_ _3918_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7002_ _3087_ _3089_ _3090_ _3091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5194_ _1265_ _1260_ _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_50_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8953_ _0026_ net11 ci_adder.instruction_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4830__A1 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7904_ _3840_ _3841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8884_ _0431_ net34 ci_adder.output_memory\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7835_ _3779_ _3784_ _3786_ _3787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_65_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6583__A1 _2694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4978_ _1122_ _1129_ _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7766_ _2471_ _3632_ _3729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6717_ _2824_ _2827_ _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7697_ ci_adder.value_i\[11\] _3629_ _3671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6648_ _2758_ _2759_ _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6579_ _2619_ _2625_ _2692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4897__A1 _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8318_ _3703_ _3524_ _4091_ _4092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9298_ _0559_ net46 ci_adder.stream_o\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9301__CLK net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7686__I1 ci_adder.uut_simple_neuron.x3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8249_ ci_adder.uut_simple_neuron.titan_id_6\[18\] _4055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_126_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5301__A2 ci_adder.uut_simple_neuron.x2\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8346__S _4070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5065__A1 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5950_ _2066_ _2072_ _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4812__A1 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4901_ _1012_ _1015_ _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5881_ _2002_ _2005_ _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_62_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7620_ ci_adder.normalised_stream_write_address\[0\] _0698_ _3602_ _3605_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4832_ _0984_ _0987_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_117_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4763_ _0886_ _0889_ _0917_ _0884_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_7551_ _3546_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6502_ _2591_ _2615_ _2616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6317__A1 _1956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4694_ _0852_ _0853_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7482_ _3479_ ci_adder.uut_simple_neuron.x0\[9\] _3475_ _3478_ _3480_ _3489_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__8306__A2 _4071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6433_ _2542_ _2547_ _2548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9221_ _0087_ net26 ci_adder.uut_simple_neuron.titan_id_2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9152_ _0244_ net76 ci_adder.uut_simple_neuron.titan_id_4\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6364_ _2145_ _2300_ _2480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6295_ _2359_ _2372_ _2412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5315_ _1427_ _1458_ _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8103_ _3945_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9083_ _0536_ net54 ci_adder.output_val_internal\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5246_ _1110_ _1343_ _1391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8034_ internal_ih.byte3\[5\] internal_ih.byte2\[5\] _3908_ _3910_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_110_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5177_ _1296_ _1323_ _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4583__I _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8936_ _0023_ net9 ci_adder.address_i\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8867_ _0414_ net50 ci_adder.output_memory\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8545__A2 _4212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8798_ _0345_ net20 internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_7818_ spi_interface_cvonk.SCLK_r\[1\] _3771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_121_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7749_ _3714_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8841__CLK net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8481__A1 _4165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8991__CLK net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5598__A2 ci_adder.uut_simple_neuron.x3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_106_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_115_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5100_ _1248_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6080_ ci_adder.uut_simple_neuron.x3\[17\] _2200_ _2201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_57_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8472__A1 ci_adder.output_val_internal\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__A1 _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5031_ ci_adder.uut_simple_neuron.x2\[18\] ci_adder.uut_simple_neuron.x2\[19\] _1181_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_57_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8076__S _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_124_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5589__A2 _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6982_ _3070_ _3071_ _3074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8721_ _0276_ net72 ci_adder.uut_simple_neuron.x3\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5933_ _2056_ _2057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_87_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5864_ _1752_ _1964_ _1988_ _1989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_91_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8652_ ci_adder.stream_o\[11\] ci_adder.output_memory\[11\] _4323_ _4325_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4815_ _0935_ _0941_ _0811_ _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout20_I net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7603_ _3589_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8583_ _4260_ _4277_ _4278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5795_ _1915_ _1921_ _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_56_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7534_ _3531_ _3529_ _3530_ _3533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4746_ ci_adder.uut_simple_neuron.x2\[6\] _0809_ _0903_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_114_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4677_ _0836_ _0837_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7465_ _3469_ _3470_ _3474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6416_ _2529_ _2498_ _2530_ _2531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9204_ _0069_ net83 ci_adder.uut_simple_neuron.titan_id_2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7396_ _3417_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8864__CLK net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6347_ _2420_ _2426_ _2463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9135_ _0169_ net91 ci_adder.uut_simple_neuron.titan_id_4\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6278_ _2347_ _2349_ _2395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9066_ _0519_ net56 ci_adder.output_val_internal\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5229_ _1372_ _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8017_ internal_ih.byte2\[5\] internal_ih.byte1\[5\] _3897_ _3901_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_123_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5202__I ci_adder.uut_simple_neuron.x2\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8919_ _0048_ net6 ci_adder.value_i\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8518__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5201__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6701__A1 ci_adder.uut_simple_neuron.x3\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5268__A1 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4600_ _0724_ ci_adder.uut_simple_neuron.x2\[5\] _0730_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_5_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5580_ _1711_ _1713_ _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5743__A2 _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7483__B _3479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ _0700_ _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4462_ internal_ih.byte1\[0\] _0648_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7250_ _3296_ _3297_ _3298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6201_ _2269_ _2268_ _2319_ _2320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_96_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7181_ _3235_ _3236_ _3239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4393_ _0619_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6132_ ci_adder.uut_simple_neuron.x3\[17\] _2251_ _2252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5259__A1 ci_adder.uut_simple_neuron.x2\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6063_ _2181_ _2183_ _2184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_84_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5014_ _0713_ _1160_ _1164_ _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_fanout68_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6965_ ci_adder.uut_simple_neuron.titan_id_4\[14\] ci_adder.uut_simple_neuron.titan_id_3\[14\]
+ _3060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5431__A1 ci_adder.uut_simple_neuron.x2\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5916_ _1774_ _2003_ _2039_ _2040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8704_ _0259_ net82 ci_adder.uut_simple_neuron.x3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_52_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6896_ ci_adder.uut_simple_neuron.titan_id_4\[3\] ci_adder.uut_simple_neuron.titan_id_3\[3\]
+ _3002_ _3003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_48_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8635_ ci_adder.stream_o\[3\] ci_adder.output_memory\[3\] _4312_ _4316_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5847_ _0163_ _1871_ _1928_ _1973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_90_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5778_ _1874_ _1888_ _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8566_ ci_adder.output_memory\[21\] _4258_ _4264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4729_ _0860_ _0863_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7517_ _3508_ ci_adder.uut_simple_neuron.x0\[15\] _3518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8497_ _0697_ _4207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_121_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7448_ ci_adder.uut_simple_neuron.x0\[3\] _3452_ _3460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7379_ ci_adder.uut_simple_neuron.titan_id_1\[23\] ci_adder.uut_simple_neuron.titan_id_0\[23\]
+ _3404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9118_ _0183_ net29 ci_adder.uut_simple_neuron.titan_id_0\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8531__S1 _4207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9049_ ci_adder.input_memory\[1\]\[17\] net38 ci_adder.uut_simple_neuron.titan_id_1\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9192__CLK net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4473__A2 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__A2 _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7478__A2 ci_adder.uut_simple_neuron.x0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6989__A1 ci_adder.uut_simple_neuron.titan_id_4\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5661__A1 _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6750_ _2860_ _2780_ _2861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5701_ _1814_ _1829_ _1813_ _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6681_ _2517_ _2707_ _2788_ _2791_ _2792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_73_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5632_ _1735_ _1737_ _1763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8420_ _3751_ ci_adder.input_memory\[1\]\[27\] _4139_ _4148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5563_ _1684_ _1693_ _1698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8351_ _4108_ _3817_ _3770_ _4109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_5_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9065__CLK net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7302_ ci_adder.uut_simple_neuron.titan_id_1\[9\] ci_adder.uut_simple_neuron.titan_id_0\[9\]
+ ci_adder.uut_simple_neuron.titan_id_1\[8\] ci_adder.uut_simple_neuron.titan_id_0\[8\]
+ _3340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4514_ ci_adder.instruction_i\[0\] ci_adder.instruction_i\[1\] _0684_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5494_ _1602_ _1633_ _1634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8282_ ci_adder.uut_simple_neuron.x0\[0\] _4072_ _4073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7233_ ci_adder.uut_simple_neuron.titan_id_2\[25\] ci_adder.uut_simple_neuron.titan_id_5\[25\]
+ _3283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4445_ _0597_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_111_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7164_ _3223_ _3224_ _3225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4376_ _0608_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6115_ _2228_ _2234_ _2235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_95_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8902__CLK net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7095_ ci_adder.uut_simple_neuron.titan_id_2\[5\] ci_adder.uut_simple_neuron.titan_id_5\[5\]
+ ci_adder.uut_simple_neuron.titan_id_2\[4\] ci_adder.uut_simple_neuron.titan_id_5\[4\]
+ _3167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6046_ _2073_ _2166_ _2167_ _2168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_107_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5404__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7997_ _3890_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6948_ _3046_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6879_ _2908_ _2915_ _2988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8618_ _0704_ _4305_ _4306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_106_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8549_ ci_adder.output_val_internal\[18\] _4249_ _4250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5643__A1 ci_adder.uut_simple_neuron.x3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_15_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5546__B _1682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7320__A1 _3354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8925__CLK net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4437__A2 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7920_ _3645_ _3841_ _3850_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8084__S _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7851_ internal_ih.spi_rx_byte_i\[6\] _3787_ _3798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6802_ _2292_ _2307_ _2912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_34_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4994_ _1109_ _1132_ _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7782_ _3741_ ci_adder.uut_simple_neuron.x3\[25\] _3692_ _3742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6733_ _1684_ _2776_ _2843_ _2844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_102_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6664_ _2773_ _2775_ _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_46_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5615_ _1728_ _1734_ _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8403_ _4116_ _4139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6595_ _2582_ _2708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_103_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5546_ _1678_ _1681_ _1682_ _1683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8334_ _3741_ ci_adder.uut_simple_neuron.x0\[25\] _4091_ _4100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5477_ _1531_ _1615_ _1616_ _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8265_ ci_adder.uut_simple_neuron.titan_id_6\[26\] _4063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7216_ _3267_ _3268_ _3269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4428_ _0639_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_113_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5873__A1 ci_adder.uut_simple_neuron.x3\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7862__A2 internal_ih.spi_rx_byte_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8196_ _3966_ _4021_ _4022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7147_ ci_adder.uut_simple_neuron.titan_id_2\[13\] ci_adder.uut_simple_neuron.titan_id_5\[13\]
+ _3211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8498__S0 _4206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4359_ internal_ih.current_instruction\[1\] internal_ih.current_instruction\[2\]
+ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8662__I1 ci_adder.output_memory\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7078_ ci_adder.uut_simple_neuron.titan_id_2\[3\] ci_adder.uut_simple_neuron.titan_id_5\[3\]
+ _3152_ _3153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5625__A1 _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6029_ _2150_ _2151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_96_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9230__CLK net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5928__A2 _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout30 net31 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout74 net75 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4600__A2 ci_adder.uut_simple_neuron.x2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout63 net69 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_12_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout41 net53 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout52 net53 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_36_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout85 net86 net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_9_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8948__CLK net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5864__A1 _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7801__S _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6216__I _2334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6380_ _1715_ _2495_ _2496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5400_ _1470_ _1541_ _1542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5331_ _1444_ _1452_ _1474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9103__CLK net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8050_ internal_ih.byte4\[5\] internal_ih.byte3\[5\] _3908_ _3918_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7001_ ci_adder.uut_simple_neuron.titan_id_4\[20\] ci_adder.uut_simple_neuron.titan_id_3\[20\]
+ _3090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5262_ _1406_ _1407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5193_ _1337_ _1338_ _1339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8952_ _0025_ net10 ci_adder.instruction_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7903_ _3839_ _3840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8883_ _0430_ net55 ci_adder.output_memory\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7834_ spi_interface_cvonk.SS_r\[1\] _3786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_93_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7765_ ci_adder.value_i\[22\] _3613_ _3727_ _3728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6716_ _2247_ _2826_ _2827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4977_ _1123_ _1128_ _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7696_ _3493_ _3663_ _3670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6647_ _2141_ _2674_ _2759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6578_ _2622_ _2624_ _2691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_115_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4897__A2 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5529_ _1666_ _1667_ _1668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8317_ _4070_ _4091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_9297_ _0558_ net46 ci_adder.stream_o\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8332__I0 _3736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8248_ _4054_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7835__A2 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8179_ _3963_ ci_adder.stream_o\[4\] ci_adder.stream_o\[20\] _3965_ _4006_ _4007_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__8635__I1 ci_adder.output_memory\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8399__I0 _3703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6023__A1 _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_25_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7771__A1 _3619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4585__A1 _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5837__A1 _1956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__A2 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5880_ _2004_ _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_88_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4900_ _1047_ _1053_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_48_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6014__A1 _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4831_ _0985_ _0944_ _0986_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7762__A1 ci_adder.uut_simple_neuron.x0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4762_ _0892_ _0916_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7550_ _3539_ ci_adder.uut_simple_neuron.x0\[21\] _3545_ _3546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_16_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6501_ _2610_ _2614_ _2615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4693_ _0850_ _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7481_ ci_adder.uut_simple_neuron.x0\[9\] _3487_ _3488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_43_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6432_ _2360_ _2477_ _2546_ _2547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9220_ _0086_ net26 ci_adder.uut_simple_neuron.titan_id_2\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9151_ _0243_ net76 ci_adder.uut_simple_neuron.titan_id_4\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6363_ _2470_ _2478_ _2479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8102_ internal_ih.byte7\[6\] internal_ih.byte6\[6\] _3825_ _3945_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6294_ _2359_ _2372_ _2411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5314_ _1430_ _1457_ _1458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9082_ _0535_ net54 ci_adder.output_val_internal\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5245_ _1110_ _1343_ _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8033_ _3909_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_110_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5176_ _1298_ _1322_ _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8935_ _0022_ net9 ci_adder.address_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8866_ _0413_ net50 ci_adder.output_memory\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7817_ spi_interface_cvonk.SS_r\[1\] _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_8797_ _0344_ net19 internal_ih.byte1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7753__A1 _3619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9149__CLK net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4567__A1 _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7748_ _3713_ _2250_ _3692_ _3714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7679_ _3612_ _3654_ _3655_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_22_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9299__CLK net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8246__I _4053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7744__A1 _3524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4558__A1 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6483__A1 _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5030_ _1157_ _1167_ _1179_ _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8472__A2 _4170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6981_ ci_adder.uut_simple_neuron.titan_id_4\[17\] ci_adder.uut_simple_neuron.titan_id_3\[17\]
+ _3073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_73_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5932_ _1803_ _2055_ _2056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8720_ _0275_ net72 ci_adder.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__8092__S _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8607__S0 _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5863_ _1754_ _1843_ _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_48_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8651_ _4324_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5794_ _1805_ _1920_ _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4814_ _0935_ _0941_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8582_ ci_adder.uut_simple_neuron.x0\[24\] ci_adder.input_memory\[1\]\[24\] ci_adder.uut_simple_neuron.x2\[24\]
+ _2538_ _4252_ _4253_ _4277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_28_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7602_ _3585_ _3588_ _3589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4745_ _0787_ ci_adder.uut_simple_neuron.x2\[8\] _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_56_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7533_ _3529_ _3530_ _3531_ _3532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_44_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout13_I internal_ih.got_all_data vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4676_ _0712_ ci_adder.uut_simple_neuron.x2\[9\] _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7464_ _3473_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8160__A1 _3966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6415_ _2462_ _2488_ _2530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9203_ _0068_ net68 ci_adder.uut_simple_neuron.titan_id_2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7395_ _3415_ _3416_ _3417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_4_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6346_ _2430_ _2434_ _2461_ _2462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9134_ _0168_ net91 ci_adder.uut_simple_neuron.titan_id_4\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9065_ _0518_ net61 ci_adder.output_val_internal\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6277_ _2338_ _2392_ _2393_ _2394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_11_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8016_ _3900_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5228_ _1034_ _1373_ _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5159_ _1224_ _1228_ _1306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_123_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8918_ _0047_ net10 ci_adder.value_i\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8849_ _0396_ net41 internal_ih.current_instruction\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4960__A1 _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8151__A1 _3966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6701__A2 ci_adder.uut_simple_neuron.x3\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8541__I3 ci_adder.uut_simple_neuron.x3\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4712__A1 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5268__A2 _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9314__CLK net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6768__A2 _2856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7764__B _3599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4530_ _0696_ _0699_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_123_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4461_ _0656_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6200_ _2265_ _2267_ _2319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_110_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4703__B2 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7180_ ci_adder.uut_simple_neuron.titan_id_2\[19\] ci_adder.uut_simple_neuron.titan_id_5\[19\]
+ _3238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6131_ _2200_ _2250_ _2251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4392_ _0601_ net14 _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_0_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5259__A2 ci_adder.uut_simple_neuron.x2\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6062_ _1675_ _2182_ _2183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_84_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5013_ _0713_ _1161_ _1163_ _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7956__A1 _3736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6964_ _3059_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5915_ _1776_ _1878_ _2039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5431__A2 ci_adder.uut_simple_neuron.x2\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8703_ _0258_ net82 ci_adder.uut_simple_neuron.x3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6895_ _2998_ _3000_ _3001_ _3002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_52_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5846_ _1906_ _1927_ _1972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8634_ _4315_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8831__CLK net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5777_ _0163_ _1871_ _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8565_ _4257_ _4259_ _4262_ _4263_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_90_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4728_ _0885_ _0886_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8496_ _0698_ _4206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7516_ ci_adder.uut_simple_neuron.x0\[15\] ci_adder.uut_simple_neuron.x0\[16\] _3517_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_114_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4659_ _0803_ _0820_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7447_ ci_adder.uut_simple_neuron.x0\[5\] _3459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_4_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7378_ _3399_ _3401_ _3402_ _3403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6329_ _2379_ _2444_ _2383_ _2445_ _2446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_9117_ _0182_ net33 ci_adder.uut_simple_neuron.titan_id_0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9048_ ci_adder.input_memory\[1\]\[16\] net37 ci_adder.uut_simple_neuron.titan_id_1\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_80_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4933__A1 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7970__I1 ci_adder.uut_simple_neuron.x2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__B2 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8854__CLK net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5700_ _1765_ _1780_ _1829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_58_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6680_ _2785_ _2789_ _2790_ _2791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6889__I _2997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5631_ _1738_ _1740_ _1760_ _1762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_73_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5562_ _1692_ _1697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__4924__A1 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8350_ spi_interface_cvonk.SS_r\[2\] _4108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7301_ _3329_ _3338_ _3339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4513_ _0683_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8281_ _4070_ _4072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5493_ _1629_ _1632_ _1633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7232_ _3269_ _3281_ _3282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4444_ _0647_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7163_ _3220_ _3221_ _3224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4375_ internal_ih.byte7\[2\] _0603_ _0607_ net14 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_fanout80_I net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6114_ _2231_ _2233_ _2234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6429__A1 _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7094_ ci_adder.uut_simple_neuron.titan_id_2\[5\] ci_adder.uut_simple_neuron.titan_id_5\[5\]
+ _3166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6045_ _2165_ _2117_ _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7996_ internal_ih.byte1\[3\] internal_ih.byte0\[3\] _3886_ _3890_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6947_ ci_adder.uut_simple_neuron.titan_id_4\[11\] ci_adder.uut_simple_neuron.titan_id_3\[11\]
+ _3045_ _3046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_64_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6878_ _2911_ _2987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5829_ _1917_ _1919_ _1955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_91_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5168__A1 ci_adder.uut_simple_neuron.x2\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8617_ ci_adder.uut_simple_neuron.x0\[31\] ci_adder.input_memory\[1\]\[31\] ci_adder.uut_simple_neuron.x2\[31\]
+ ci_adder.uut_simple_neuron.x3\[31\] _0698_ _0697_ _4305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_36_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4915__A1 _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8548_ _4161_ _4249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_118_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8479_ ci_adder.output_memory\[6\] _4163_ _4192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5340__A1 _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8877__CLK net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5634__A2 _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7850_ internal_ih.spi_tx_byte_o\[5\] _3779_ _3784_ internal_ih.spi_rx_byte_i\[5\]
+ _3797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6801_ _2909_ _2910_ _2911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_34_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4993_ _1144_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7709__S _3632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9032__CLK net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7781_ _3738_ _3740_ _3741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6732_ _2773_ _2775_ _2843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_102_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7139__A2 ci_adder.uut_simple_neuron.titan_id_5\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6663_ _1792_ _2774_ _2775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_85_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9182__CLK net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5614_ _1728_ _1734_ _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6898__A1 ci_adder.uut_simple_neuron.titan_id_4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7934__I1 ci_adder.uut_simple_neuron.x2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8402_ _4138_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6594_ _2576_ _2644_ _2707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5545_ _1678_ _1680_ _1682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_53_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8333_ _4099_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5476_ _0711_ ci_adder.uut_simple_neuron.x2\[29\] _1616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7847__B1 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8264_ _4062_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7215_ ci_adder.uut_simple_neuron.titan_id_2\[25\] ci_adder.uut_simple_neuron.titan_id_5\[25\]
+ _3268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4427_ internal_ih.byte5\[7\] _0635_ _0632_ internal_ih.byte1\[7\] _0639_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8195_ _3962_ ci_adder.stream_o\[14\] _4021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_113_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5873__A2 ci_adder.uut_simple_neuron.x3\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7146_ ci_adder.uut_simple_neuron.titan_id_2\[13\] ci_adder.uut_simple_neuron.titan_id_5\[13\]
+ _3210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8498__S1 _4207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4358_ internal_ih.current_instruction\[0\] internal_ih.current_instruction\[1\]
+ internal_ih.current_instruction\[2\] _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_7077_ _3148_ _3150_ _3151_ _3152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5625__A2 _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6028_ _1878_ _2149_ _2150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__A1 ci_adder.uut_simple_neuron.x2\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7979_ internal_ih.byte0\[3\] internal_ih.spi_rx_byte_i\[3\] _3877_ _3881_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_83_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout31 net40 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout20 net21 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout64 net69 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_12_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout42 net53 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout53 net92 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_37_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout86 net89 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout75 net80 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_12_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__A1 _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7838__B1 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5552__A1 _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5330_ _1471_ _1472_ _1473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5261_ _1401_ _1402_ _1405_ _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_50_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7000_ ci_adder.uut_simple_neuron.titan_id_4\[20\] ci_adder.uut_simple_neuron.titan_id_3\[20\]
+ _3089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5192_ _1318_ _1320_ _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8951_ _0016_ net8 ci_adder.address_i\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7902_ _3610_ _3838_ _3839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8882_ _0429_ net54 ci_adder.output_memory\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8557__A1 _4211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7833_ internal_ih.spi_tx_byte_o\[0\] _3779_ _3784_ internal_ih.spi_rx_byte_i\[0\]
+ _3785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_fanout43_I net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7764_ _3725_ _3726_ _3599_ _3727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6715_ _2254_ _2825_ _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4976_ _1126_ _1127_ _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_63_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5791__A1 ci_adder.uut_simple_neuron.x3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7695_ ci_adder.uut_simple_neuron.x0\[10\] _3657_ ci_adder.uut_simple_neuron.x0\[11\]
+ _3669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6646_ _2147_ _2673_ _2758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6577_ _1726_ _1728_ _2635_ _2690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_116_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7682__B ci_adder.uut_simple_neuron.x0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_115_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5528_ _1481_ _1624_ _1667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8316_ _4090_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9296_ _0557_ net48 ci_adder.stream_o\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5459_ _1597_ _1598_ _1599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8247_ ci_adder.uut_simple_neuron.titan_id_6\[17\] _4054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8178_ _3966_ _4005_ _4006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7129_ ci_adder.uut_simple_neuron.titan_id_2\[10\] ci_adder.uut_simple_neuron.titan_id_5\[10\]
+ _3197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_126_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8915__CLK net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4585__A2 ci_adder.uut_simple_neuron.x2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8200__C _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5837__A2 _1962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8539__A1 _4211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4830_ _0870_ _0945_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4761_ _0918_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6500_ _2094_ _2613_ _2614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4692_ ci_adder.uut_simple_neuron.x2\[9\] ci_adder.uut_simple_neuron.x2\[10\] _0852_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_56_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7514__A2 ci_adder.uut_simple_neuron.x0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7480_ ci_adder.uut_simple_neuron.x0\[10\] _3487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_15_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6431_ _2545_ _2476_ _2546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9150_ _0242_ net78 ci_adder.uut_simple_neuron.titan_id_4\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6362_ _2360_ _2477_ _2478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5313_ _1433_ _1456_ _1457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8101_ _3944_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6293_ _2403_ _2409_ _2410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_12_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9081_ _0534_ net54 ci_adder.output_val_internal\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5244_ _1387_ _1388_ _1389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8032_ internal_ih.byte3\[4\] internal_ih.byte2\[4\] _3908_ _3909_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_110_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5175_ _1301_ _1321_ _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6846__B ci_adder.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8617__I2 ci_adder.uut_simple_neuron.x2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8934_ _0021_ net9 ci_adder.address_i\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8938__CLK net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8865_ _0412_ net51 ci_adder.output_memory\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7816_ _3769_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8796_ _0343_ net20 internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_121_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ _1085_ _1110_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7747_ _3710_ _3711_ _3712_ _3713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7678_ ci_adder.uut_simple_neuron.x3\[8\] _3617_ _3655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8002__I0 internal_ih.byte1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6629_ _2739_ _2666_ _2740_ _2741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_62_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6600__I _2712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9279_ _0144_ net33 ci_adder.uut_simple_neuron.titan_id_6\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5755__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4558__A2 _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7807__S _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9243__CLK net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6180__A1 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6483__A2 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7680__A1 _3479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4494__A1 internal_ih.byte2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6980_ _3072_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8480__I0 _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5931_ _1805_ _1917_ _2055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_73_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8607__S1 _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5862_ _1952_ _1968_ _1986_ _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8650_ ci_adder.stream_o\[10\] ci_adder.output_memory\[10\] _4323_ _4324_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5793_ _1917_ _1919_ _1920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4813_ _0808_ _0965_ _0968_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8581_ ci_adder.output_memory\[24\] _4258_ _4276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_38_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7601_ _3582_ _3586_ _3587_ _3581_ _3588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4744_ _0901_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_60_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7532_ ci_adder.uut_simple_neuron.x0\[17\] ci_adder.uut_simple_neuron.x0\[18\] _3531_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_126_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4675_ _0815_ _0835_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9202_ _0067_ net85 ci_adder.uut_simple_neuron.titan_id_2\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7463_ _3469_ _3470_ _3472_ _3473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_31_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6414_ _2462_ _2488_ _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7394_ ci_adder.uut_simple_neuron.titan_id_1\[26\] ci_adder.uut_simple_neuron.titan_id_0\[26\]
+ _3416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6345_ _2417_ _2429_ _2461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9133_ _0167_ net87 ci_adder.uut_simple_neuron.titan_id_4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6276_ _2341_ _2375_ _2393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_47_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_9064_ _0517_ net61 ci_adder.output_val_internal\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5227_ _1370_ _1199_ _1372_ _1373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7671__A1 _3608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8015_ internal_ih.byte2\[4\] internal_ih.byte1\[4\] _3897_ _3900_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_71_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8760__CLK net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4485__A1 internal_ih.byte2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5158_ _1224_ _1228_ _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_47_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5089_ _1119_ _1219_ _1237_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_123_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9116__CLK net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8917_ _0046_ net6 ci_adder.value_i\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_56_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8848_ _0395_ net19 internal_ih.current_instruction\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8779_ _0326_ net28 ci_adder.uut_simple_neuron.x2\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_65_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7662__A1 ci_adder.uut_simple_neuron.x3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5976__A1 _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8142__A2 _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ internal_ih.byte0\[7\] _0648_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4391_ _0618_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6130_ ci_adder.uut_simple_neuron.x3\[19\] _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_21_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6061_ _1792_ _1810_ _2182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9139__CLK net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9203__D _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__A1 internal_ih.byte1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7653__A1 _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5012_ _1162_ _1160_ _1163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7956__A2 _3846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5967__A1 _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6963_ _3057_ _3058_ _3059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9289__CLK net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5914_ _1991_ _2036_ _2037_ _2038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6894_ ci_adder.uut_simple_neuron.titan_id_4\[2\] ci_adder.uut_simple_neuron.titan_id_3\[2\]
+ _3001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8702_ _0257_ net58 ci_adder.uut_simple_neuron.x3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_52_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5845_ _1945_ _1970_ _1971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_105_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5719__A1 _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8633_ ci_adder.stream_o\[2\] ci_adder.output_memory\[2\] _4312_ _4315_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8381__A2 _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5776_ _1896_ _1856_ _1895_ _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8564_ ci_adder.output_val_internal\[20\] _4249_ _4263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4727_ _0869_ _0871_ _0883_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7515_ _3516_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8133__A2 _3964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8495_ ci_adder.output_memory\[9\] _4163_ _4205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4658_ _0804_ _0819_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7446_ _3458_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7892__A1 _3826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4589_ _0747_ _0753_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9116_ _0181_ net36 ci_adder.uut_simple_neuron.titan_id_0\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7377_ ci_adder.uut_simple_neuron.titan_id_1\[22\] ci_adder.uut_simple_neuron.titan_id_0\[22\]
+ _3402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8516__S0 _4206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6328_ _2386_ _2445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6259_ _2278_ _2312_ _2377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7644__A1 _3612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9047_ ci_adder.input_memory\[1\]\[15\] net37 ci_adder.uut_simple_neuron.titan_id_1\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4458__A1 internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__A1 _1723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4630__A1 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_73_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6374__A1 _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5630_ _1761_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5561_ _1686_ _1687_ _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7066__I _3143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5492_ _1630_ _1631_ _1632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7300_ _3330_ _3335_ _3338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8115__A2 _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4512_ ci_adder.uut_simple_neuron.x0\[0\] ci_adder.uut_simple_neuron.x0\[1\] _0683_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8280_ _4070_ _4071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_124_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7231_ _3275_ _3277_ _3281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8098__S _3825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4443_ internal_ih.byte6\[7\] _0602_ _0619_ internal_ih.byte2\[7\] _0647_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_111_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7162_ ci_adder.uut_simple_neuron.titan_id_2\[16\] ci_adder.uut_simple_neuron.titan_id_5\[16\]
+ _3223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4374_ internal_ih.byte4\[2\] internal_ih.byte3\[2\] _0599_ _0607_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6429__A2 _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6113_ _0162_ _2232_ _2233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7093_ _3157_ _3158_ _3163_ _3165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6044_ _2165_ _2117_ _2166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout73_I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7995_ _3889_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _3035_ _3041_ _3044_ _3045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_76_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7685__B _3660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6877_ _2984_ _2985_ _2986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5828_ _1922_ _1924_ _1953_ _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_64_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8616_ ci_adder.output_memory\[31\] _0703_ _4304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5759_ _1886_ _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8547_ _4214_ _4247_ _4248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_118_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8106__A2 _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6668__A2 _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7865__A1 internal_ih.spi_rx_byte_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9304__CLK net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8478_ _4162_ _4188_ _4190_ _4191_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7429_ _3445_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__A1 _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8593__A2 _4285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6356__A1 _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6108__A1 _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7815__S _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6659__A2 _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7856__A1 internal_ih.spi_rx_byte_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7084__A2 ci_adder.uut_simple_neuron.titan_id_5\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8408__I0 _3723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6800_ _2247_ _2826_ _2910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8971__CLK net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4992_ _1138_ _1143_ _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7780_ ci_adder.uut_simple_neuron.x0\[25\] _3730_ _3739_ _3614_ _3740_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_34_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6731_ _2801_ _2841_ _2842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_102_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6662_ _1801_ _1810_ _2774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5613_ _1722_ _1743_ _1744_ _1745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8401_ _3708_ ci_adder.input_memory\[1\]\[18\] _4122_ _4138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6593_ _2646_ _2705_ _2706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_73_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8332_ _3736_ ci_adder.uut_simple_neuron.x0\[24\] _4091_ _4099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5544_ _1675_ _1680_ _1681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_30_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5475_ _0711_ ci_adder.uut_simple_neuron.x2\[29\] _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8263_ ci_adder.uut_simple_neuron.titan_id_6\[25\] _4062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7214_ ci_adder.uut_simple_neuron.titan_id_2\[25\] ci_adder.uut_simple_neuron.titan_id_5\[25\]
+ _3267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4426_ _0638_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8194_ _3979_ _4019_ _4020_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7145_ _3209_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_113_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4357_ internal_ih.current_instruction\[5\] internal_ih.current_instruction\[4\]
+ internal_ih.current_instruction\[7\] internal_ih.current_instruction\[6\] _0592_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__5086__A1 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7076_ ci_adder.uut_simple_neuron.titan_id_2\[2\] ci_adder.uut_simple_neuron.titan_id_5\[2\]
+ _3151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6027_ _1880_ _1997_ _2149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6822__A2 _2931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7978_ _3804_ _3877_ _3880_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6929_ _3018_ _3021_ _3030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout21 net24 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout10 net11 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_119_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout65 net66 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_49_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout54 net57 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_12_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout43 net44 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout32 net39 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_37_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout76 net80 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout87 net88 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_92_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7838__B2 internal_ih.spi_rx_byte_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6510__A1 _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8844__CLK net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5077__A1 ci_adder.uut_simple_neuron.x2\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8994__CLK net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5001__A1 _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5552__A2 _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5260_ _0712_ _1403_ _1404_ _1349_ _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_23_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_10_Left_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5191_ _1309_ _1336_ _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8950_ _0015_ net8 ci_adder.address_i\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7901_ _3608_ _3605_ _3603_ _3838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8881_ _0428_ net82 ci_adder.output_memory\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7832_ _3783_ _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4975_ _0718_ ci_adder.uut_simple_neuron.x2\[18\] _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout36_I net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7763_ ci_adder.uut_simple_neuron.x0\[22\] _3721_ _3726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6714_ _2364_ _2745_ _2744_ _2825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_74_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5791__A2 ci_adder.uut_simple_neuron.x3\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7694_ _3617_ _3667_ _3668_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6645_ _2755_ _2756_ _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6576_ _2652_ _2688_ _2689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6740__A1 _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5543__A2 _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8867__CLK net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5527_ _1479_ _1623_ _1666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8315_ _3697_ ci_adder.uut_simple_neuron.x0\[16\] _4076_ _4090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9295_ _0556_ net48 ci_adder.stream_o\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8246_ _4053_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5458_ _1470_ _1582_ _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5389_ ci_adder.uut_simple_neuron.x2\[27\] ci_adder.uut_simple_neuron.x2\[28\] _1531_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4409_ internal_ih.byte4\[7\] _0623_ _0620_ internal_ih.byte0\[7\] _0629_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8177_ _3962_ ci_adder.stream_o\[12\] _4005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7128_ _3190_ _3191_ _3192_ _3194_ _3195_ _3196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_7059_ _3138_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_126_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5231__A1 _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4585__A3 ci_adder.uut_simple_neuron.x2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8484__A1 ci_adder.output_memory\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5298__A1 ci_adder.uut_simple_neuron.x2\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9022__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9172__CLK net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5470__A1 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7211__A2 ci_adder.uut_simple_neuron.titan_id_5\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4760_ _0891_ _0917_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6970__A1 ci_adder.uut_simple_neuron.titan_id_4\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4691_ _0718_ ci_adder.uut_simple_neuron.x2\[9\] _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8011__I1 internal_ih.byte1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _2467_ _2543_ _2544_ _2545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6361_ _2473_ _2476_ _2477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5312_ _1437_ _1455_ _1456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8100_ internal_ih.byte7\[5\] internal_ih.byte6\[5\] _3825_ _3944_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6292_ _2406_ _2408_ _2409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9080_ _0533_ net56 ci_adder.output_val_internal\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5243_ _1335_ _1362_ _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8031_ _3818_ _3908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_110_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5174_ _1318_ _1320_ _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5461__A1 _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8933_ _0020_ net9 ci_adder.address_i\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8864_ _0411_ net49 ci_adder.output_memory\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7815_ _3768_ ci_adder.uut_simple_neuron.x3\[31\] _3611_ _3769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8795_ _0342_ net20 internal_ih.byte1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_121_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4958_ _0811_ _1083_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_46_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7746_ ci_adder.value_i\[19\] _3659_ _3712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4889_ _0714_ _1042_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7677_ ci_adder.value_i\[8\] _3613_ _3653_ _3654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__8002__I1 internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6628_ _2662_ _2667_ _2740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9045__CLK net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6559_ _2656_ _2671_ _2672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7913__S _3846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8466__A1 _4165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9278_ _0143_ net32 ci_adder.uut_simple_neuron.titan_id_6\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8229_ ci_adder.uut_simple_neuron.titan_id_6\[8\] _4045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8069__I1 internal_ih.byte4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_2_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A2 _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_123_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6180__A2 _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7680__A2 ci_adder.uut_simple_neuron.x0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8654__S _4323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7807__I1 ci_adder.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5930_ _2047_ _2053_ _2054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ _1954_ _1967_ _1986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7600_ ci_adder.uut_simple_neuron.x0\[28\] ci_adder.uut_simple_neuron.x0\[29\] _3587_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_118_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5792_ ci_adder.uut_simple_neuron.x3\[10\] _1918_ _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_4
X_4812_ _0939_ _0967_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8580_ _4257_ _4272_ _4274_ _4275_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_83_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4743_ _0899_ _0900_ _0895_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_60_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7531_ ci_adder.uut_simple_neuron.x0\[15\] _3524_ ci_adder.uut_simple_neuron.x0\[16\]
+ _3530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7462_ _3459_ _3469_ _3471_ _3472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6413_ _2526_ _2527_ _2528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4674_ _0709_ _0790_ _0834_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_71_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9201_ _0095_ net68 ci_adder.uut_simple_neuron.titan_id_2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7393_ _3411_ _3412_ _3414_ _3415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6344_ _2410_ _2436_ _2459_ _2460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9132_ _0166_ net91 ci_adder.uut_simple_neuron.titan_id_4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6275_ _2341_ _2375_ _2392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8905__CLK net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8628__I _3601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9063_ _0516_ net48 ci_adder.output_val_internal\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5226_ _1198_ _1245_ _1371_ _1372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8014_ _3899_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_71_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4485__A2 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5157_ _1265_ _1302_ _1303_ _1304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_79_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5088_ _1223_ _1232_ _1236_ _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8620__A1 _4170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8916_ _0045_ net6 ci_adder.value_i\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8363__I _4116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8847_ _0394_ net41 internal_ih.current_instruction\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8778_ _0325_ net72 ci_adder.uut_simple_neuron.x2\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_19_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7729_ _3697_ _2098_ _3692_ _3698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__I2 ci_adder.uut_simple_neuron.x2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8439__A1 _3966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5673__A1 ci_adder.uut_simple_neuron.x3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7662__A2 _3617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5897__I _2021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5425__A1 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5976__A2 _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9210__CLK net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8470__S0 _4166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7973__I0 internal_ih.byte0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8928__CLK net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7780__C _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ internal_ih.byte7\[7\] _0603_ _0617_ net14 _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8448__I _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6060_ _2179_ _2180_ _2181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4467__A2 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5011_ ci_adder.uut_simple_neuron.x2\[18\] ci_adder.uut_simple_neuron.x2\[19\] _1162_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6962_ ci_adder.uut_simple_neuron.titan_id_4\[14\] ci_adder.uut_simple_neuron.titan_id_3\[14\]
+ _3058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5913_ _1993_ _2006_ _2037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8701_ _0256_ net82 ci_adder.uut_simple_neuron.x3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6893_ ci_adder.uut_simple_neuron.titan_id_4\[2\] ci_adder.uut_simple_neuron.titan_id_3\[2\]
+ _3000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_52_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5844_ _1947_ _1969_ _1970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_105_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5719__A2 _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8632_ _4314_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7964__I0 _3757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8563_ _4260_ _4261_ _4262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5775_ _1863_ _1899_ _1901_ _1902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7514_ _3508_ ci_adder.uut_simple_neuron.x0\[15\] _3515_ _3516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_44_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4726_ _0884_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8494_ _4162_ _4200_ _4202_ _4204_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4657_ _0805_ _0818_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7445_ _3453_ _3457_ _3458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7376_ ci_adder.uut_simple_neuron.titan_id_1\[22\] ci_adder.uut_simple_neuron.titan_id_0\[22\]
+ _3401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_2_Left_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6327_ _2380_ _2318_ _2444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4588_ _0709_ _0749_ _0752_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__8516__S1 _4207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9115_ _0180_ net36 ci_adder.uut_simple_neuron.titan_id_0\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6258_ _2338_ _2341_ _2375_ _2376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7644__A2 _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9046_ ci_adder.input_memory\[1\]\[14\] net60 ci_adder.uut_simple_neuron.titan_id_1\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _2307_ _2308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5209_ _1353_ _1354_ _1355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5958__A2 _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6080__A1 ci_adder.uut_simple_neuron.x3\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4394__B2 internal_ih.byte0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8683__I1 ci_adder.output_memory\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__A1 _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7946__I0 _3713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8750__CLK net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ _1686_ _1687_ _1694_ _1695_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_81_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5491_ _1560_ _1580_ _1631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4511_ _0682_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8371__I0 _3631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4442_ _0646_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7230_ _3280_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5885__A1 _1945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7161_ _3222_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4373_ _0606_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6112_ _1836_ _1851_ _2232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_95_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7092_ _3164_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6043_ _2116_ _2165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9256__CLK net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout66_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7994_ internal_ih.byte1\[2\] internal_ih.byte0\[2\] _3886_ _3889_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_37_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _3042_ _3043_ _3044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6876_ _2921_ _2932_ _2985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_66_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5827_ _1915_ _1921_ _1953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8615_ _4170_ _4300_ _4302_ _4303_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_36_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5758_ _1884_ _1885_ _1886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_8546_ ci_adder.uut_simple_neuron.x0\[18\] ci_adder.input_memory\[1\]\[18\] ci_adder.uut_simple_neuron.x2\[18\]
+ _2200_ _4206_ _4207_ _4247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_118_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4709_ _0868_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8477_ ci_adder.output_val_internal\[5\] _4170_ _4191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5689_ _1781_ _1784_ _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_32_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7428_ ci_adder.uut_simple_neuron.titan_id_1\[31\] ci_adder.uut_simple_neuron.titan_id_0\[31\]
+ _3444_ _3445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5876__A1 _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7359_ _3387_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9029_ _0512_ net41 internal_ih.expected_byte_count\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8290__A2 _4071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4851__A2 ci_adder.uut_simple_neuron.x2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6053__A1 _1723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4603__A2 ci_adder.uut_simple_neuron.x2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6356__A2 _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9129__CLK net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4367__A1 internal_ih.current_instruction\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5867__A1 _1956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8656__I1 ci_adder.output_memory\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5619__A1 ci_adder.uut_simple_neuron.x3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8662__S _4323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6730_ _2830_ _2840_ _2841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4991_ _1141_ _1142_ _1143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_86_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6661_ _1677_ _1700_ _2771_ _2772_ _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_102_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6592_ _2701_ _2704_ _2705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5612_ _1735_ _1737_ _1744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8400_ _4137_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5543_ ci_adder.uut_simple_neuron.x3\[1\] _1679_ _1680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8331_ _4098_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5858__A1 _1721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5474_ _1613_ _1614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8262_ _4061_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4425_ internal_ih.byte5\[6\] _0635_ _0632_ internal_ih.byte1\[6\] _0638_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8193_ internal_ih.spi_tx_byte_o\[5\] _3978_ _4020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7213_ _3266_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_92_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7144_ ci_adder.uut_simple_neuron.titan_id_2\[13\] ci_adder.uut_simple_neuron.titan_id_5\[13\]
+ _3208_ _3209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4356_ _0591_ internal_ih.got_all_data vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4530__A1 _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8647__I1 ci_adder.output_memory\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5086__A2 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7075_ ci_adder.uut_simple_neuron.titan_id_2\[2\] ci_adder.uut_simple_neuron.titan_id_5\[2\]
+ _3150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6026_ _2141_ _2147_ _2148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5060__I _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6586__A2 _2698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7977_ internal_ih.byte0\[2\] _3877_ _3880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6928_ _3029_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout11 internal_ih.got_all_data net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout22 net24 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_107_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6859_ _2966_ _2967_ _2968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout55 net57 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout33 net39 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout44 net53 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout77 net80 net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout88 net89 net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout66 net69 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_12_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8529_ _4211_ _4230_ _4232_ _4233_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_103_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7651__S _3632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6274__A1 _1682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8281__I _4070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4588__A1 _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8326__I0 _3723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4512__A1 ci_adder.uut_simple_neuron.x0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _1314_ _1317_ _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7900_ _3826_ _3837_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_92_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8880_ _0427_ net56 ci_adder.output_memory\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7831_ _3780_ _3782_ _3783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4974_ _1095_ _1125_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7762_ ci_adder.uut_simple_neuron.x0\[22\] _3721_ _3725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6713_ _2823_ _2824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7693_ ci_adder.uut_simple_neuron.x3\[10\] _3632_ _3668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout29_I net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6644_ _1778_ _2684_ _2756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_63_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7736__S _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8190__A1 _3811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6575_ _2677_ _2687_ _2688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5526_ _1614_ _1617_ _1664_ _1665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8314_ _4089_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9294_ _0555_ net48 ci_adder.stream_o\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5457_ _1556_ _1581_ _1597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8245_ ci_adder.uut_simple_neuron.titan_id_6\[16\] _4053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4408_ _0628_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8493__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5388_ ci_adder.uut_simple_neuron.x2\[28\] _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_8176_ _3979_ _4003_ _4004_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_74_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7127_ ci_adder.uut_simple_neuron.titan_id_2\[9\] ci_adder.uut_simple_neuron.titan_id_5\[9\]
+ _3195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7058_ ci_adder.uut_simple_neuron.titan_id_4\[30\] ci_adder.uut_simple_neuron.titan_id_3\[30\]
+ _3137_ _3138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_6009_ _2092_ _2107_ _2131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_126_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7508__A1 ci_adder.uut_simple_neuron.x0\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4990__A1 _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8811__CLK net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8181__A1 _3811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4742__A1 _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5298__A2 ci_adder.uut_simple_neuron.x2\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8961__CLK net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7113__C ci_adder.uut_simple_neuron.titan_id_5\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9317__CLK net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8209__C _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5470__A2 ci_adder.uut_simple_neuron.x2\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4690_ ci_adder.uut_simple_neuron.x2\[9\] ci_adder.uut_simple_neuron.x2\[10\] _0850_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8172__A1 _3811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8562__I3 ci_adder.uut_simple_neuron.x3\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6360_ _2365_ _2475_ _2476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5311_ _1441_ _1454_ _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6291_ _1704_ _2407_ _2408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6486__A1 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8387__S _4122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8030_ _3907_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5242_ _1339_ _1361_ _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_110_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5173_ _1119_ _1319_ _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_46_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6238__A1 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 spi_clock_i net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8932_ _0019_ net9 ci_adder.address_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8863_ _0410_ net46 internal_ih.spi_tx_byte_o\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7814_ ci_adder.value_i\[31\] _3767_ _3614_ _3768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6410__A1 _2491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8834__CLK net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8794_ _0341_ net22 internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_121_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4957_ _1076_ _1099_ _1108_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7745_ _3536_ _3700_ _3614_ _3711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4888_ _1017_ _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4972__A1 _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7676_ _3613_ _3652_ _3653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_22_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6627_ _2664_ _2739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6558_ _2669_ _2670_ _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7910__A1 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6489_ _2424_ _2602_ _2603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5509_ _1611_ _1619_ _1648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9277_ _0142_ net33 ci_adder.uut_simple_neuron.titan_id_6\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8228_ _4044_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8159_ _3962_ ci_adder.stream_o\[10\] _3989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7977__A1 internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5204__A2 ci_adder.uut_simple_neuron.x2\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7901__A1 _3608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8457__A2 _4170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8480__I2 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8857__CLK net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5860_ _1678_ _1984_ _1985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4811_ _0909_ _0966_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7196__A2 ci_adder.uut_simple_neuron.titan_id_5\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5791_ ci_adder.uut_simple_neuron.x3\[11\] ci_adder.uut_simple_neuron.x3\[12\] _1918_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_7_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4742_ _0899_ _0894_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_60_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7530_ ci_adder.uut_simple_neuron.x0\[16\] _3524_ _3519_ _3521_ _3517_ _3529_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_7_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4673_ ci_adder.uut_simple_neuron.x2\[6\] _0787_ ci_adder.uut_simple_neuron.x2\[8\]
+ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7461_ _3465_ _3466_ _3464_ _3471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_126_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6412_ _1725_ _1728_ _2456_ _2527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_114_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9200_ _0094_ net67 ci_adder.uut_simple_neuron.titan_id_2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7392_ ci_adder.uut_simple_neuron.titan_id_1\[25\] ci_adder.uut_simple_neuron.titan_id_0\[25\]
+ _3414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6343_ _2413_ _2435_ _2459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9131_ _0165_ net87 ci_adder.uut_simple_neuron.titan_id_4\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6274_ _1682_ _2337_ _2391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9062_ _0515_ net45 internal_ih.data_pointer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5225_ _1285_ _1325_ _1371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8013_ internal_ih.byte2\[3\] internal_ih.byte1\[3\] _3897_ _3899_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_71_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5156_ _1016_ _1091_ _1259_ _1303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5087_ _1222_ _1234_ _1235_ _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_27_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8915_ _0043_ net10 ci_adder.value_i\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_123_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8846_ _0393_ net15 internal_ih.byte7\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5989_ _2111_ _2112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_109_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5198__A1 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8777_ _0324_ net72 ci_adder.uut_simple_neuron.x2\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__9012__CLK net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7728_ _3619_ _3694_ _3695_ _3696_ _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__8136__A1 _3966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__I3 ci_adder.uut_simple_neuron.x3\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6698__A1 ci_adder.uut_simple_neuron.x3\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9127__D ci_adder.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7659_ _3452_ _3627_ _3459_ _3639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_62_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6870__A1 _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8611__A2 _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5425__A2 ci_adder.uut_simple_neuron.x2\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5189__A1 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8470__S1 _4167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4936__A1 _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7973__I1 internal_ih.spi_rx_byte_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7102__A2 ci_adder.uut_simple_neuron.titan_id_5\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5010_ ci_adder.uut_simple_neuron.x2\[18\] _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5664__A2 _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6861__A1 _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6961_ _3053_ _3055_ _3056_ _3057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_88_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8700_ _0255_ net82 ci_adder.uut_simple_neuron.x3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__9035__CLK net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5912_ _1993_ _2006_ _2036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6892_ _2999_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_52_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5843_ _1952_ _1968_ _1969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_105_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8631_ ci_adder.stream_o\[1\] ci_adder.output_memory\[1\] _4312_ _4314_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__9185__CLK net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4927__A1 _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7964__I1 _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8562_ _3539_ ci_adder.input_memory\[1\]\[20\] ci_adder.uut_simple_neuron.x2\[20\]
+ ci_adder.uut_simple_neuron.x3\[20\] _4252_ _4253_ _4261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5774_ _1865_ _1898_ _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7513_ _3509_ _3512_ _3514_ _3515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout11_I internal_ih.got_all_data vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4725_ _0869_ _0871_ _0883_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8493_ ci_adder.output_val_internal\[8\] _4203_ _4204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4656_ _0793_ _0802_ _0817_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_25_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7444_ _3454_ _3455_ _3456_ _3457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_114_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4587_ _0750_ _0751_ _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7375_ _3400_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6326_ _2321_ _2383_ _2443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9114_ _0179_ net38 ci_adder.uut_simple_neuron.titan_id_0\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5104__A1 _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6257_ _2351_ _2374_ _2375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9045_ ci_adder.input_memory\[1\]\[13\] net60 ci_adder.uut_simple_neuron.titan_id_1\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6188_ _1997_ _2306_ _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6852__A1 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5208_ ci_adder.uut_simple_neuron.x2\[23\] _1185_ _1267_ _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_4_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5139_ _1243_ _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6080__A2 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8829_ _0376_ net15 internal_ih.byte5\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4918__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4394__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_112_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_95_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9058__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_121_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8596__A1 ci_adder.output_memory\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6532__I _2645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7946__I1 ci_adder.uut_simple_neuron.x2\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7628__I _3599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5582__A1 _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ _1562_ _1579_ _1630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4510_ internal_ih.byte3\[7\] _0597_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4441_ internal_ih.byte6\[6\] _0602_ _0619_ internal_ih.byte2\[6\] _0646_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8520__A1 ci_adder.output_memory\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7160_ _3220_ _3221_ _3222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6111_ _2229_ _2230_ _2231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4372_ internal_ih.byte7\[1\] _0603_ _0605_ net14 _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_95_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8395__S _4122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7091_ _3162_ _3163_ _3164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6042_ _2160_ _2163_ _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5637__A2 _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_107_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout59_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7993_ _3888_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6944_ ci_adder.uut_simple_neuron.titan_id_4\[10\] ci_adder.uut_simple_neuron.titan_id_3\[10\]
+ ci_adder.uut_simple_neuron.titan_id_4\[9\] ci_adder.uut_simple_neuron.titan_id_3\[9\]
+ _3043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_88_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6875_ _2924_ _2931_ _2984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_66_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8614_ ci_adder.output_val_internal\[30\] _4161_ _4303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5826_ _1699_ _1951_ _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5757_ _1713_ _1774_ _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8545_ ci_adder.output_memory\[18\] _4212_ _4246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4708_ _0864_ _0867_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_45_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8198__S0 _3964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8476_ _4165_ _4189_ _4190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_118_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5688_ _1781_ _1784_ _1818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5325__A1 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7427_ _3440_ _3441_ _3443_ _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_102_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4639_ _0761_ _0798_ _0799_ _0781_ _0800_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_4_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7358_ _3385_ _3386_ _3387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6309_ _2252_ _2425_ _2426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9200__CLK net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7289_ _3325_ _3326_ _3327_ _3328_ _3329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_9028_ _0511_ net18 ci_adder.input_memory\[1\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__A3 ci_adder.uut_simple_neuron.x2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6053__A2 _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8918__CLK net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7250__A1 _3296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8050__I0 internal_ih.byte4\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8189__S0 _3964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5316__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7856__A3 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5867__A2 _1962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6816__A1 _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5619__A2 ci_adder.uut_simple_neuron.x3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6292__A2 _2408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4990_ _1034_ _1068_ _1103_ _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_86_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6660_ _1770_ _1772_ _2772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_102_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6591_ _2583_ _2702_ _2703_ _2704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5611_ _1735_ _1737_ _1743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5555__A1 _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4358__A2 internal_ih.current_instruction\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5542_ ci_adder.uut_simple_neuron.x3\[2\] _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_53_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8330_ _3733_ ci_adder.uut_simple_neuron.x0\[23\] _4091_ _4098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5473_ _1612_ _1530_ ci_adder.uut_simple_neuron.x2\[30\] _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__9223__CLK net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9225__D _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8261_ ci_adder.uut_simple_neuron.titan_id_6\[24\] _4061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7212_ _3264_ _3265_ _3266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4424_ _0637_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8192_ ci_adder.stream_o\[29\] _3959_ _4018_ _4019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7143_ _3204_ _3205_ _3207_ _3208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4355_ _0583_ internal_ih.received_byte_count\[2\] _0585_ _0590_ _0591_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_113_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7074_ _3149_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6025_ _1999_ _2146_ _2147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_68_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7976_ _3879_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6927_ _3027_ _3028_ _3029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xfanout12 internal_ih.got_all_data net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6858_ _2905_ _2916_ _2967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout56 net57 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout23 net24 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout45 net47 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout34 net39 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout78 net79 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5809_ _1866_ _1934_ _1935_ _1936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5546__A1 _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout89 net90 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout67 net69 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_9_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6789_ _2886_ _2898_ _2899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8528_ ci_adder.output_val_internal\[14\] _4203_ _4233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7932__S _3855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8459_ ci_adder.output_memory\[2\] _4163_ _4176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7471__A1 _3470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6026__A2 _2147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5785__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8023__I0 internal_ih.byte3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9246__CLK net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8582__S0 _4252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7462__A1 _3459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7830_ spi_interface_cvonk.state\[2\] _3781_ _3782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_47_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7765__A2 _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4973_ _1016_ _1124_ _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7761_ _3724_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6712_ _2806_ _2822_ _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7692_ ci_adder.value_i\[10\] _3613_ _3666_ _3667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_19_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6643_ _2135_ _2150_ _2755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7517__A2 ci_adder.uut_simple_neuron.x0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6574_ _2680_ _2686_ _2687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_6_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8140__C _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5525_ _1573_ _1618_ _1664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8313_ _3691_ ci_adder.uut_simple_neuron.x0\[15\] _4076_ _4089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9293_ _0554_ net46 ci_adder.stream_o\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5456_ _1595_ _1596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8244_ _4052_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4407_ internal_ih.byte4\[6\] _0623_ _0620_ internal_ih.byte0\[6\] _0628_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5387_ _1487_ _1488_ _1529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8175_ internal_ih.spi_tx_byte_o\[3\] _3978_ _4004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_74_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7126_ _3180_ _3181_ _3193_ _3194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_10_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7057_ _3133_ _3135_ _3136_ _3137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7453__A1 _3459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6008_ _2080_ _2129_ _2130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9119__CLK net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7959_ _3870_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4415__I _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7692__A1 ci_adder.value_i\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6183__A1 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8786__CLK net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8668__S _4323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6290_ _1950_ _1965_ _2407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5310_ _1400_ _1453_ _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6486__A2 ci_adder.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5241_ _0994_ _1364_ _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_110_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5172_ _0808_ _1083_ _1304_ _1319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xinput2 spi_cs_i net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8931_ _0018_ net9 ci_adder.address_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8862_ _0409_ net44 internal_ih.spi_tx_byte_o\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7738__A2 _3629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5749__A1 ci_adder.uut_simple_neuron.x3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout41_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8793_ _0340_ net20 internal_ih.byte1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7813_ ci_adder.uut_simple_neuron.x0\[31\] _3593_ _3760_ _3767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7744_ _3524_ _3695_ ci_adder.uut_simple_neuron.x0\[19\] _3710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4956_ _1078_ _1098_ _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4421__B2 internal_ih.byte1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4887_ _1003_ _1010_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4972__A2 ci_adder.uut_simple_neuron.x2\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7675_ _3479_ _3647_ _3652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6626_ _2540_ _2737_ _2738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6174__A1 _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6557_ _2300_ _2302_ _2473_ _2670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7910__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5508_ _1620_ _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8546__S0 _4206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6488_ _2599_ _2601_ _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9276_ _0141_ net32 ci_adder.uut_simple_neuron.titan_id_6\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _1562_ _1579_ _1580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7674__A1 _3612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4488__A1 internal_ih.byte2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8227_ ci_adder.uut_simple_neuron.titan_id_6\[7\] _4044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8158_ _3979_ _3987_ _3988_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7109_ _3158_ _3163_ _3179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8089_ _3938_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_87_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A2 ci_adder.uut_simple_neuron.x2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7665__A1 _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4479__A1 internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7191__I _3247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8465__I0 ci_adder.uut_simple_neuron.x0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__A1 _1960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8480__I3 ci_adder.uut_simple_neuron.x3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4810_ _0874_ _0931_ _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5790_ ci_adder.uut_simple_neuron.x3\[9\] _1879_ _1916_ _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_68_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4403__B2 internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4403__A1 internal_ih.byte4\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4741_ ci_adder.uut_simple_neuron.x2\[12\] _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_60_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4672_ _0714_ _0810_ _0816_ _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_56_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7460_ ci_adder.uut_simple_neuron.x0\[7\] _3470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_44_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6411_ _2524_ _2525_ _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9130_ _0164_ net87 ci_adder.uut_simple_neuron.titan_id_4\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7391_ _3413_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6342_ _2454_ _2457_ _2458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6273_ _2381_ _2379_ _2389_ _2390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7656__A1 ci_adder.uut_simple_neuron.x3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9061_ ci_adder.input_memory\[1\]\[29\] net25 ci_adder.uut_simple_neuron.titan_id_1\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5224_ _1068_ _1103_ _1370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8012_ _3898_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout89_I net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5155_ _1225_ _1261_ _1055_ _1302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5086_ _0712_ _1233_ _1221_ _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_16_Left_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8801__CLK net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8914_ _0042_ net10 ci_adder.value_i\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_123_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4642__A1 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8845_ _0392_ net15 internal_ih.byte7\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8951__CLK net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5988_ _2033_ _2076_ _2110_ _2111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5198__A2 _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8776_ _0323_ net72 ci_adder.uut_simple_neuron.x2\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_47_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4939_ _1055_ _1057_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7727_ ci_adder.value_i\[16\] _3659_ _3696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7658_ _3452_ _3459_ _3627_ _3638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__9307__CLK net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_25_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6609_ _2689_ _2721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6698__A2 ci_adder.uut_simple_neuron.x3\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7895__A1 _3826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7589_ ci_adder.uut_simple_neuron.x0\[26\] ci_adder.uut_simple_neuron.x0\[27\] _3578_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_15_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9259_ _0154_ net51 ci_adder.uut_simple_neuron.titan_id_6\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7940__S _3855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5425__A3 _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8375__A2 _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4936__A2 ci_adder.uut_simple_neuron.x2\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_43_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8011__S _3897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7638__A1 _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8824__CLK net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6310__A1 _2100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6613__A2 _2687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6960_ ci_adder.uut_simple_neuron.titan_id_4\[13\] ci_adder.uut_simple_neuron.titan_id_3\[13\]
+ _3056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5911_ _2033_ _2034_ _2035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6891_ ci_adder.uut_simple_neuron.titan_id_4\[2\] ci_adder.uut_simple_neuron.titan_id_3\[2\]
+ _2998_ _2999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_49_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8366__A2 _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5842_ _1954_ _1967_ _1968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6377__A1 _1956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8630_ _4313_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5773_ _1900_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8561_ _0704_ _4260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_118_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6129__A1 _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4724_ _0845_ _0882_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7512_ _3502_ _3508_ _3514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8492_ _4161_ _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4655_ _0810_ _0816_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7443_ ci_adder.uut_simple_neuron.x0\[1\] ci_adder.uut_simple_neuron.x0\[2\] _3456_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4586_ _0722_ ci_adder.uut_simple_neuron.x2\[4\] ci_adder.uut_simple_neuron.x2\[5\]
+ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7374_ ci_adder.uut_simple_neuron.titan_id_1\[22\] ci_adder.uut_simple_neuron.titan_id_0\[22\]
+ _3399_ _3400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_6325_ _2390_ _2441_ _2442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9113_ _0178_ net37 ci_adder.uut_simple_neuron.titan_id_0\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8677__I0 ci_adder.stream_o\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7760__S _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9044_ ci_adder.input_memory\[1\]\[12\] net60 ci_adder.uut_simple_neuron.titan_id_1\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6301__A1 _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6256_ _2353_ _2373_ _2374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6187_ _1999_ _2143_ _2306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5207_ _1221_ _1352_ _1353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_4_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5138_ _1198_ _1245_ _1286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5069_ _1055_ _1124_ _1181_ _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_94_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6368__A1 _2100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8828_ _0375_ net15 internal_ih.byte5\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8759_ _0306_ net82 ci_adder.uut_simple_neuron.x2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_63_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8293__A1 _3459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4854__A1 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4606__A1 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6359__A1 _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5031__A1 ci_adder.uut_simple_neuron.x2\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5582__A2 _1715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4440_ _0645_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8520__A2 _4212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6110_ _1801_ _2191_ _2230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4371_ internal_ih.byte4\[1\] internal_ih.byte3\[1\] _0599_ _0605_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7087__A2 ci_adder.uut_simple_neuron.titan_id_5\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7090_ ci_adder.uut_simple_neuron.titan_id_2\[5\] ci_adder.uut_simple_neuron.titan_id_5\[5\]
+ _3163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6041_ _2074_ _2161_ _2162_ _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9002__CLK net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6598__A1 _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9152__CLK net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7992_ internal_ih.byte1\[1\] internal_ih.byte0\[1\] _3886_ _3888_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6943_ ci_adder.uut_simple_neuron.titan_id_4\[10\] ci_adder.uut_simple_neuron.titan_id_3\[10\]
+ _3042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6874_ _2965_ _2968_ _2982_ _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_88_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5825_ _1704_ _1950_ _1951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8613_ _0704_ _4301_ _4302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_119_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5756_ _1711_ _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8544_ _4211_ _4242_ _4244_ _4245_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_115_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5687_ _1764_ _1817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4707_ _0865_ _0866_ _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8475_ _3459_ ci_adder.input_memory\[1\]\[5\] ci_adder.uut_simple_neuron.x2\[5\]
+ ci_adder.uut_simple_neuron.x3\[5\] _4166_ _4167_ _4189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_118_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4638_ _0783_ _0796_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7426_ ci_adder.uut_simple_neuron.titan_id_1\[30\] ci_adder.uut_simple_neuron.titan_id_0\[30\]
+ _3443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4569_ _0715_ _0722_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7357_ ci_adder.uut_simple_neuron.titan_id_1\[19\] ci_adder.uut_simple_neuron.titan_id_0\[19\]
+ _3386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6308_ _2422_ _2424_ _2425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5089__A1 _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7288_ ci_adder.uut_simple_neuron.titan_id_1\[7\] ci_adder.uut_simple_neuron.titan_id_0\[7\]
+ _3328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6239_ _1915_ _2356_ _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9027_ _0510_ net25 ci_adder.input_memory\[1\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8578__A2 _4273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5013__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9025__CLK net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9175__CLK net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6590_ _2586_ _2639_ _2703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5610_ _1738_ _1740_ _1742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5555__A2 ci_adder.uut_simple_neuron.x3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8592__I2 ci_adder.uut_simple_neuron.x2\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ ci_adder.uut_simple_neuron.x3\[0\] _1676_ _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_54_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_42_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8260_ _4060_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5472_ ci_adder.uut_simple_neuron.x2\[27\] _1612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7211_ ci_adder.uut_simple_neuron.titan_id_2\[24\] ci_adder.uut_simple_neuron.titan_id_5\[24\]
+ _3265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_30_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4423_ internal_ih.byte5\[5\] _0635_ _0632_ internal_ih.byte1\[5\] _0637_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8191_ _3960_ _4015_ _4017_ _3815_ _4018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_111_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7142_ ci_adder.uut_simple_neuron.titan_id_2\[12\] ci_adder.uut_simple_neuron.titan_id_5\[12\]
+ _3207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4354_ _0586_ _0588_ _0589_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_113_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7073_ ci_adder.uut_simple_neuron.titan_id_2\[2\] ci_adder.uut_simple_neuron.titan_id_5\[2\]
+ _3148_ _3149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6024_ _2143_ _2145_ _2146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9241__D _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout71_I net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7975_ internal_ih.byte0\[1\] internal_ih.spi_rx_byte_i\[1\] _3877_ _3879_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6926_ ci_adder.uut_simple_neuron.titan_id_4\[8\] ci_adder.uut_simple_neuron.titan_id_3\[8\]
+ _3028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6991__A1 ci_adder.uut_simple_neuron.titan_id_4\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout13 internal_ih.got_all_data net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6857_ _2883_ _2904_ _2966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout35 net39 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8032__I1 internal_ih.byte2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout24 net40 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout46 net47 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout79 net80 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5808_ _1891_ _1894_ _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6743__A1 _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6788_ _2896_ _2897_ _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout68 net69 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout57 net70 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5739_ _0162_ _1836_ _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9048__CLK net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8527_ _4214_ _4231_ _4232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8458_ _4162_ _4172_ _4174_ _4175_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_33_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7409_ _3427_ _3428_ _3429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8389_ _3677_ ci_adder.input_memory\[1\]\[12\] _4122_ _4132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9198__CLK net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4809__A1 _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5482__A1 ci_adder.uut_simple_neuron.x2\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7471__A2 _3479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5785__A2 _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8023__I1 internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7782__I0 _3741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8582__S1 _4253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7462__A2 _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8411__A1 _3728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4972_ _1011_ ci_adder.uut_simple_neuron.x2\[16\] ci_adder.uut_simple_neuron.x2\[17\]
+ _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7760_ _3723_ _2365_ _3692_ _3724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6711_ _2817_ _2821_ _2822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7691_ _3614_ _3665_ _3666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6642_ _2728_ _2753_ _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_63_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6573_ _2683_ _2685_ _2686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8312_ _4088_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5524_ _0994_ _1662_ _1663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9292_ _0553_ net48 ci_adder.stream_o\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5455_ _1593_ _1594_ _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8243_ ci_adder.uut_simple_neuron.titan_id_6\[15\] _4052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8908__CLK net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4406_ _0627_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8174_ ci_adder.stream_o\[27\] _3959_ _4002_ _4003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5386_ _1526_ _1527_ _1528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7125_ _3176_ _3183_ _3193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_74_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7056_ ci_adder.uut_simple_neuron.titan_id_4\[29\] ci_adder.uut_simple_neuron.titan_id_3\[29\]
+ _3136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_66_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6007_ _2125_ _2128_ _2129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_126_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7958_ _3741_ ci_adder.uut_simple_neuron.x2\[25\] _3840_ _3870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6909_ ci_adder.uut_simple_neuron.titan_id_4\[5\] ci_adder.uut_simple_neuron.titan_id_3\[5\]
+ _3013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7889_ internal_ih.received_byte_count\[3\] _3829_ _3831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_108_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8104__S _3825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8469__A1 ci_adder.output_memory\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7692__A2 _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9213__CLK net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5240_ _1332_ _1363_ _1385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5171_ _1309_ _1314_ _1317_ _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8930_ _0017_ net10 ci_adder.address_i\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput3 spi_pico_i net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8861_ _0408_ net42 internal_ih.spi_tx_byte_o\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5749__A2 ci_adder.uut_simple_neuron.x3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8792_ _0339_ net20 internal_ih.byte1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7994__I0 internal_ih.byte1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7812_ _3766_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4955_ _1107_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7743_ _3709_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout34_I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4421__A2 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4886_ _1039_ _1010_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7674_ _3612_ _3650_ _3651_ _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_22_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6625_ _2734_ _2736_ _2737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_116_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6556_ _2661_ _2668_ _2669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_89_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5507_ _1644_ _1645_ _1646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_76_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8546__S1 _4207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9275_ _0140_ net35 ci_adder.uut_simple_neuron.titan_id_6\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6487_ _2474_ _2600_ _2601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_14_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8226_ _4043_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5438_ _1525_ _1578_ _1579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8880__CLK net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5369_ _1500_ _1502_ _1504_ _1511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8157_ internal_ih.spi_tx_byte_o\[1\] _3979_ _3988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8088_ internal_ih.byte6\[7\] internal_ih.byte5\[7\] _3930_ _3938_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7108_ _3152_ _3155_ _3177_ _3178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7039_ _3121_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9236__CLK net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_98_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7938__S _3855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7985__I0 internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_98_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4479__A2 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5720__I _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_57_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8753__CLK net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4403__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7647__I _3608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4740_ _0811_ _0897_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4671_ _0788_ _0831_ _0815_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_126_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6410_ _2491_ _2497_ _2525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7390_ _3411_ _3412_ _3413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9109__CLK net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6341_ _1686_ _1709_ _2456_ _2457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_114_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8153__I0 ci_adder.output_val_internal\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6272_ _2376_ _2378_ _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_110_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7656__A2 _3617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9060_ ci_adder.input_memory\[1\]\[28\] net27 ci_adder.uut_simple_neuron.titan_id_1\[30\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5667__A1 _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5223_ _1367_ _1368_ _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8011_ internal_ih.byte2\[2\] internal_ih.byte1\[2\] _3897_ _3898_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5154_ _1299_ _1273_ _1300_ _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5419__A1 _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5085_ _1233_ _1221_ _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_27_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8913_ _0041_ net10 ci_adder.value_i\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_123_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8844_ _0391_ net17 internal_ih.byte7\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5987_ _2083_ _2109_ _2110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_94_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8775_ _0322_ net72 ci_adder.uut_simple_neuron.x2\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_4938_ _1089_ _1090_ _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7726_ ci_adder.uut_simple_neuron.x0\[16\] _3689_ _3695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_19_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4869_ _1000_ _1023_ _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_82_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7657_ _3612_ _3636_ _3637_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6608_ _2690_ _2697_ _2719_ _2720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7588_ ci_adder.uut_simple_neuron.x0\[26\] ci_adder.uut_simple_neuron.x0\[27\] _3577_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6539_ _2616_ _2626_ _2651_ _2652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9258_ _0153_ net63 ci_adder.uut_simple_neuron.titan_id_6\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9189_ _0222_ net76 ci_adder.uut_simple_neuron.titan_id_3\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8209_ _3960_ _4031_ _4033_ _3815_ _4034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_7_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6083__A1 _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8776__CLK net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8455__S0 _4166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7958__I0 _3741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8207__S0 _3964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7638__A2 _3617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6310__A2 _2249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__A1 _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5910_ _1725_ _2030_ _2031_ _2034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_88_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6890_ ci_adder.uut_simple_neuron.titan_id_4\[1\] ci_adder.uut_simple_neuron.titan_id_3\[1\]
+ _2998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5841_ _1963_ _1966_ _1967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5772_ _1863_ _1899_ _1900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8560_ ci_adder.output_memory\[20\] _4258_ _4259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4723_ _0872_ _0881_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7511_ _3513_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8491_ _4165_ _4201_ _4202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_32_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7442_ ci_adder.uut_simple_neuron.x0\[0\] ci_adder.uut_simple_neuron.x0\[1\] ci_adder.uut_simple_neuron.x0\[2\]
+ _3455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4654_ _0788_ _0811_ _0815_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7877__A2 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4585_ _0722_ ci_adder.uut_simple_neuron.x2\[4\] ci_adder.uut_simple_neuron.x2\[5\]
+ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_7373_ _3395_ _3396_ _3398_ _3399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9081__CLK net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6324_ _2391_ _2440_ _2441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_101_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4560__A1 _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9112_ _0177_ net38 ci_adder.uut_simple_neuron.titan_id_0\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6255_ _2357_ _2359_ _2372_ _2373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_9043_ ci_adder.input_memory\[1\]\[11\] net59 ci_adder.uut_simple_neuron.titan_id_1\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5206_ ci_adder.uut_simple_neuron.x2\[23\] _1267_ _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6186_ _2298_ _2304_ _2305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5137_ _1281_ _1284_ _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_4_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8799__CLK net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5068_ _1215_ _1189_ _1216_ _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_84_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6368__A2 _2249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7565__A1 ci_adder.uut_simple_neuron.x0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8827_ _0374_ net15 internal_ih.byte5\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8758_ _0305_ net58 ci_adder.uut_simple_neuron.x2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7709_ _3680_ ci_adder.uut_simple_neuron.x3\[13\] _3632_ _3681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_124_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8689_ ci_adder.stream_o\[29\] ci_adder.output_memory\[29\] _4334_ _4344_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4551__A1 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8293__A2 _4072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6359__A2 _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5031__A2 ci_adder.uut_simple_neuron.x2\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4370_ _0604_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8941__CLK net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8284__A2 _4072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6040_ _2112_ _2114_ _2162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7991_ _3887_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6942_ _3036_ _3039_ _3041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_37_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6873_ _2737_ _2971_ _2981_ _2982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5824_ _1732_ _1803_ _1949_ _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_76_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_17_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8612_ ci_adder.uut_simple_neuron.x0\[30\] ci_adder.input_memory\[1\]\[30\] ci_adder.uut_simple_neuron.x2\[30\]
+ ci_adder.uut_simple_neuron.x3\[30\] _0698_ _0697_ _4301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_91_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5755_ _1876_ _1882_ _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_56_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8543_ ci_adder.output_val_internal\[17\] _4203_ _4245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5686_ _1813_ _1815_ _1816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4706_ _0801_ _0821_ _0827_ _0842_ _0823_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_8474_ ci_adder.output_memory\[5\] _4163_ _4188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4637_ _0783_ _0796_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_62_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7425_ _3442_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4568_ _0727_ _0733_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7356_ _3383_ _3384_ _3385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6307_ ci_adder.uut_simple_neuron.x3\[20\] _2423_ _2424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7287_ ci_adder.uut_simple_neuron.titan_id_1\[7\] ci_adder.uut_simple_neuron.titan_id_0\[7\]
+ ci_adder.uut_simple_neuron.titan_id_1\[6\] ci_adder.uut_simple_neuron.titan_id_0\[6\]
+ _3327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4499_ _0676_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6238_ _1921_ _2355_ _2356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_9026_ _0509_ net25 ci_adder.input_memory\[1\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6169_ _2281_ _2287_ _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_90_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_71_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7946__S _3855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8338__I0 _3751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6513__A2 _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8964__CLK net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8017__S _3897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8592__I3 ci_adder.uut_simple_neuron.x3\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5540_ _1677_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_54_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5471_ _1609_ _1610_ _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7210_ ci_adder.uut_simple_neuron.titan_id_2\[23\] ci_adder.uut_simple_neuron.titan_id_5\[23\]
+ _3253_ _3261_ _3263_ _3264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4422_ _0636_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_112_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8190_ _3811_ _4016_ _4017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7141_ _3206_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4353_ internal_ih.expected_byte_count\[3\] _0584_ internal_ih.received_byte_count\[5\]
+ internal_ih.received_byte_count\[1\] _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_39_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7072_ _3144_ _3145_ _3147_ _3148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6023_ _2050_ _2144_ _2145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4818__A2 ci_adder.uut_simple_neuron.x2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout64_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7974_ _3878_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6925_ _3025_ _3026_ _3027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8837__CLK net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6856_ _2963_ _2964_ _2965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout36 net38 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout47 net53 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout25 net27 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_119_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5807_ _1891_ _1894_ _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6787_ _2473_ _2476_ _2664_ _2897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xfanout58 net70 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout69 net70 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8987__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5738_ _1814_ _1829_ _1813_ _1856_ _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8526_ _3508_ ci_adder.input_memory\[1\]\[14\] ci_adder.uut_simple_neuron.x2\[14\]
+ ci_adder.uut_simple_neuron.x3\[14\] _4206_ _4207_ _4231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_45_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5669_ _1796_ _1797_ _1798_ _1799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_103_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8457_ ci_adder.output_val_internal\[1\] _4170_ _4175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8388_ _4131_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7408_ ci_adder.uut_simple_neuron.titan_id_1\[28\] ci_adder.uut_simple_neuron.titan_id_0\[28\]
+ _3428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7339_ _3366_ _3368_ _3370_ _3371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9009_ _0492_ net60 ci_adder.input_memory\[1\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5482__A2 _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7759__A1 _3619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4365__S _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_109_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__A1 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7782__I1 ci_adder.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8487__A2 _4170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9142__CLK net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_118_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5473__A2 _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8411__A2 _4117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6422__A1 _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4971_ _0713_ _1096_ _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6710_ _2422_ _2820_ _2821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7690_ _3663_ _3664_ _3665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6641_ _2731_ _2747_ _2752_ _2753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_73_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6572_ _1778_ _2684_ _2685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8311_ _3685_ _3508_ _4076_ _4088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5523_ _1643_ _1646_ _1661_ _1662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_6_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9291_ _0552_ net49 ci_adder.stream_o\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5454_ _0994_ _1584_ _1594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8242_ _4051_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5385_ _1482_ _1490_ _1527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5161__A1 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4405_ internal_ih.byte4\[5\] _0623_ _0620_ internal_ih.byte0\[5\] _0627_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8173_ _3960_ _3999_ _4001_ _3815_ _4002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_112_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9252__D _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7124_ _3185_ _3188_ _3192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_74_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7055_ ci_adder.uut_simple_neuron.titan_id_4\[29\] ci_adder.uut_simple_neuron.titan_id_3\[29\]
+ _3135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6006_ _2127_ _2128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6464__I _2578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7957_ _1348_ _3841_ _3869_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9015__CLK net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4975__A1 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6908_ _3012_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7888_ internal_ih.received_byte_count\[3\] _3829_ _3830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_119_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6839_ _2349_ _2372_ _2948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9165__CLK net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8509_ _4211_ _4213_ _4216_ _4217_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_21_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5391__A1 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5170_ _1308_ _1316_ _1317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_110_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput4 sys_clock_i net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9038__CLK net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8860_ _0407_ net42 internal_ih.spi_tx_byte_o\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8791_ _0338_ net20 internal_ih.byte1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7811_ _3765_ ci_adder.uut_simple_neuron.x3\[30\] _3611_ _3766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__9188__CLK net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4954_ _1103_ _1106_ _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7742_ _3708_ _2200_ _3692_ _3709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7994__I1 internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout27_I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4885_ _0811_ _1037_ _1038_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9247__D _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7673_ ci_adder.uut_simple_neuron.x3\[7\] _3617_ _3651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4532__I _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6624_ ci_adder.uut_simple_neuron.x3\[25\] _2735_ _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6555_ _2662_ _2667_ _2668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5382__A1 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5506_ _0994_ _1635_ _1645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_76_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9274_ _0139_ net35 ci_adder.uut_simple_neuron.titan_id_6\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6486_ _2538_ ci_adder.uut_simple_neuron.x3\[25\] _2600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7123__A2 ci_adder.uut_simple_neuron.titan_id_5\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8225_ ci_adder.uut_simple_neuron.titan_id_6\[6\] _4043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5437_ _1565_ _1577_ _1578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5368_ _1500_ _1502_ _1510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8156_ ci_adder.stream_o\[25\] _3959_ _3986_ _3987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5299_ _1442_ _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8087_ _3937_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7107_ ci_adder.uut_simple_neuron.titan_id_2\[3\] ci_adder.uut_simple_neuron.titan_id_5\[3\]
+ _3177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7038_ _3119_ _3120_ _3121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6634__A1 _2364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8989_ _0472_ net27 ci_adder.uut_simple_neuron.x0\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_93_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8139__A1 _3811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7954__S _3840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5125__A1 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8614__A2 _4161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8465__I2 _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8378__A1 _3645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4939__A1 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8025__S _3897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4670_ _0808_ _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_56_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8550__A1 _4211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6340_ _1686_ _2455_ _2456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6271_ _2388_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_122_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5667__A2 _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6864__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5222_ _1329_ _1330_ _1365_ _1368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8010_ _3825_ _3897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_110_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5153_ _1274_ _1277_ _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_71_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5084_ ci_adder.uut_simple_neuron.x2\[21\] _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8912_ _0040_ net10 ci_adder.value_i\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8369__A1 _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8843_ _0390_ net16 internal_ih.byte7\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_27_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5986_ _2085_ _2108_ _2109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_93_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8774_ _0321_ net29 ci_adder.uut_simple_neuron.x2\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_47_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4937_ _1011_ ci_adder.uut_simple_neuron.x2\[16\] ci_adder.uut_simple_neuron.x2\[17\]
+ _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_47_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7725_ ci_adder.uut_simple_neuron.x0\[16\] _3689_ _3694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4868_ _1019_ _1022_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_82_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7656_ ci_adder.uut_simple_neuron.x3\[4\] _3617_ _3637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ _2693_ _2696_ _2719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4799_ _0831_ _0911_ _0954_ _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_7587_ ci_adder.uut_simple_neuron.x0\[27\] ci_adder.uut_simple_neuron.x0\[28\] _3576_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6538_ _2591_ _2615_ _2651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6469_ _2526_ _2527_ _2583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9257_ _0152_ net51 ci_adder.uut_simple_neuron.titan_id_6\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9188_ _0221_ net76 ci_adder.uut_simple_neuron.titan_id_3\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8208_ _3811_ _4032_ _4033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_7_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8139_ _3811_ _3970_ _3971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7958__I1 ci_adder.uut_simple_neuron.x2\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8455__S1 _4167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5594__A1 _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8383__I1 ci_adder.input_memory\[1\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8720__CLK net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5840_ _1965_ _1966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8870__CLK net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5771_ _1865_ _1898_ _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5585__A1 _1699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4722_ _0879_ _0880_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8490_ _3479_ ci_adder.input_memory\[1\]\[8\] ci_adder.uut_simple_neuron.x2\[8\]
+ ci_adder.uut_simple_neuron.x3\[8\] _4166_ _4167_ _4201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7510_ _3509_ _3512_ _3513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7441_ ci_adder.uut_simple_neuron.x0\[3\] _3454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_126_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4653_ _0812_ _0813_ _0814_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_72_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4584_ _0748_ _0730_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7372_ ci_adder.uut_simple_neuron.titan_id_1\[21\] ci_adder.uut_simple_neuron.titan_id_0\[21\]
+ _3398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6323_ _2394_ _2439_ _2440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9111_ _0176_ net37 ci_adder.uut_simple_neuron.titan_id_0\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6254_ _2362_ _2369_ _2371_ _2372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_9042_ ci_adder.input_memory\[1\]\[10\] net59 ci_adder.uut_simple_neuron.titan_id_1\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ _1349_ _1350_ _1351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6185_ _2195_ _2303_ _2304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_5136_ _1282_ _1283_ _1284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5067_ _1182_ _1188_ _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_84_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8826_ _0373_ net17 internal_ih.byte5\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5969_ _2054_ _2057_ _2091_ _2092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_94_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5576__A1 ci_adder.uut_simple_neuron.x3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8757_ _0304_ net83 ci_adder.uut_simple_neuron.x2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_51_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7708_ ci_adder.value_i\[13\] _3679_ _3614_ _3680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8688_ _4343_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8514__A1 _4211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7639_ _3612_ _3621_ _3622_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4551__A2 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9309_ _0570_ net45 ci_adder.stream_o\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8743__CLK net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7253__A1 _3296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8053__I0 internal_ih.byte4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5567__A1 _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9249__CLK net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6819__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7492__A1 ci_adder.uut_simple_neuron.x0\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7795__A2 _3612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7990_ internal_ih.byte1\[0\] internal_ih.byte0\[0\] _3886_ _3887_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6941_ _3040_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6872_ _2974_ _2977_ _2980_ _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_88_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5823_ _1948_ _1923_ _1949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8611_ ci_adder.output_memory\[30\] _0703_ _4300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8542_ _4214_ _4243_ _4244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5754_ _1776_ _1881_ _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_91_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5685_ _1765_ _1780_ _1814_ _1815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4705_ _0827_ _0842_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8473_ _4162_ _4184_ _4186_ _4187_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4636_ _0766_ _0787_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4540__I ci_adder.uut_simple_neuron.x2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7424_ _3440_ _3441_ _3442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8766__CLK net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7355_ _3380_ _3381_ _3384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6306_ ci_adder.uut_simple_neuron.x3\[21\] ci_adder.uut_simple_neuron.x3\[22\] _2423_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4567_ _0709_ _0729_ _0732_ _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7286_ _3317_ _3322_ _3326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4498_ internal_ih.byte3\[1\] _0670_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6237_ _1997_ _2306_ _2354_ _2355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7483__A1 _3470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9025_ _0508_ net27 ci_adder.input_memory\[1\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6168_ _2284_ _2286_ _2287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_90_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ ci_adder.uut_simple_neuron.x2\[21\] ci_adder.uut_simple_neuron.x2\[22\] _1267_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_6099_ _2219_ _2160_ _2164_ _2168_ _2220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__7786__A2 _3608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5549__A1 _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8809_ _0356_ net23 internal_ih.byte3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5721__A1 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9071__CLK net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4460__A1 internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5470_ _0712_ ci_adder.uut_simple_neuron.x2\[29\] _1531_ _1610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_26_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4421_ internal_ih.byte5\[4\] _0635_ _0632_ internal_ih.byte1\[4\] _0636_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7701__A2 _3659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7140_ _3204_ _3205_ _3206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4352_ internal_ih.expected_byte_count\[0\] _0587_ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6287__I _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7465__A1 _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7071_ ci_adder.uut_simple_neuron.titan_id_2\[1\] ci_adder.uut_simple_neuron.titan_id_5\[1\]
+ _3147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6022_ _2098_ ci_adder.uut_simple_neuron.x3\[17\] _2144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4818__A3 ci_adder.uut_simple_neuron.x2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout57_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7973_ internal_ih.byte0\[0\] internal_ih.spi_rx_byte_i\[0\] _3877_ _3878_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6924_ _3022_ _3023_ _3026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6855_ _2298_ _2902_ _2964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout37 net38 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout15 net16 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_18_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout26 net27 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5806_ _1929_ _1932_ _1933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6786_ _2889_ _2895_ _2896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout59 net70 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout48 net49 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5737_ _1827_ _1864_ _1865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8525_ ci_adder.output_memory\[14\] _4212_ _4230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7782__S _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8456_ _4165_ _4173_ _4174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5668_ _1772_ _1778_ _1798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_79_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7407_ _3415_ _3423_ _3426_ _3427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5599_ ci_adder.uut_simple_neuron.x3\[4\] _1731_ _1732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_4
X_4619_ _0761_ _0779_ _0781_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8387_ _3672_ ci_adder.input_memory\[1\]\[11\] _4122_ _4131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_92_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7338_ ci_adder.uut_simple_neuron.titan_id_1\[15\] ci_adder.uut_simple_neuron.titan_id_0\[15\]
+ _3370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7269_ ci_adder.uut_simple_neuron.titan_id_1\[5\] ci_adder.uut_simple_neuron.titan_id_0\[5\]
+ _3311_ _3312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_9008_ _0491_ net60 ci_adder.input_memory\[1\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9094__CLK net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4445__I _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8008__I0 internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4745__A2 ci_adder.uut_simple_neuron.x2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8567__S0 _4252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4681__A1 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5473__A3 ci_adder.uut_simple_neuron.x2\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _1119_ _1121_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6640_ _2197_ _2751_ _2752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_86_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6571_ _2135_ _2150_ _2684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4736__A2 ci_adder.uut_simple_neuron.x2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7922__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5522_ _1649_ _1660_ _1661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8310_ _4087_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9290_ _0551_ net49 ci_adder.stream_o\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5453_ _1553_ _1583_ _1593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8497__I _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8241_ ci_adder.uut_simple_neuron.titan_id_6\[14\] _4051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5384_ _1483_ _1489_ _1526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4404_ _0626_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8172_ _3811_ _4000_ _4001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7123_ ci_adder.uut_simple_neuron.titan_id_2\[9\] ci_adder.uut_simple_neuron.titan_id_5\[9\]
+ _3191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_74_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7054_ _3134_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6110__A1 _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8804__CLK net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6005_ _1765_ _1770_ _2126_ _2127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6661__A2 _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4672__A1 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6413__A2 _2527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8954__CLK net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7956_ _3736_ _3846_ _3869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6907_ _3010_ _3011_ _3012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4975__A2 ci_adder.uut_simple_neuron.x2\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7887_ _3826_ _3828_ _3829_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_108_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6838_ _1915_ _2943_ _2946_ _2947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_92_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5924__A1 ci_adder.uut_simple_neuron.x3\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6769_ _2878_ _2879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8508_ ci_adder.output_val_internal\[10\] _4203_ _4217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8401__S _4122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7677__A1 ci_adder.value_i\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8439_ _3966_ _3974_ _4159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8401__I0 _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5391__A2 _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8311__S _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7668__A1 _3612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6340__A1 _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8827__CLK net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7840__A1 _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7810_ ci_adder.value_i\[30\] _3764_ _3614_ _3765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8790_ _0337_ net41 internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4953_ _1104_ _1105_ _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7741_ _3705_ _3707_ _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_47_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7672_ ci_adder.value_i\[7\] _3619_ _3649_ _3650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6623_ ci_adder.uut_simple_neuron.x3\[26\] ci_adder.uut_simple_neuron.x3\[27\] _2735_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4884_ _0965_ _0968_ _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5906__A1 _1715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ _2664_ _2666_ _2667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6485_ _2471_ _2597_ _2598_ _2599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5505_ _1599_ _1634_ _1644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9273_ _0137_ net35 ci_adder.uut_simple_neuron.titan_id_6\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7659__A1 _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5436_ _1482_ _1576_ _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_76_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8224_ _4042_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5367_ _1366_ _1418_ _1419_ _1507_ _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4893__A1 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8155_ _3960_ _3983_ _3985_ _3815_ _3986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5298_ ci_adder.uut_simple_neuron.x2\[24\] ci_adder.uut_simple_neuron.x2\[25\] _1442_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7106_ ci_adder.uut_simple_neuron.titan_id_2\[7\] ci_adder.uut_simple_neuron.titan_id_5\[7\]
+ _3176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8086_ internal_ih.byte6\[6\] internal_ih.byte5\[6\] _3930_ _3937_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7037_ ci_adder.uut_simple_neuron.titan_id_4\[27\] ci_adder.uut_simple_neuron.titan_id_3\[27\]
+ _3120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4645__A1 _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9132__CLK net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8988_ _0471_ net28 ci_adder.uut_simple_neuron.x0\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_2_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7939_ _3860_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5070__A1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7970__S _3840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6873__A2 _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8465__I3 ci_adder.uut_simple_neuron.x3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7822__A1 _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4636__A1 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8378__A2 _4117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8622__I0 _4166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6561__A1 _2147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6270_ _2383_ _2387_ _2388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5221_ _1366_ _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5152_ _1258_ _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6616__A2 _2675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9155__CLK net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5083_ _1229_ _1231_ _1232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8911_ _0039_ net12 ci_adder.value_i\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8369__A2 _4117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8842_ _0389_ net17 internal_ih.byte7\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8773_ _0320_ net73 ci_adder.uut_simple_neuron.x2\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_63_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5985_ _2089_ _2092_ _2107_ _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5052__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__I _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7724_ _3693_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4936_ _1011_ ci_adder.uut_simple_neuron.x2\[16\] ci_adder.uut_simple_neuron.x2\[17\]
+ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_117_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4867_ _1020_ _1021_ _0980_ _0978_ _0932_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XTAP_TAPCELL_ROW_82_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7655_ _3613_ _3634_ _3635_ _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6606_ _2701_ _2704_ _2718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6552__A1 ci_adder.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7586_ _3575_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6537_ _2628_ _2638_ _2649_ _2650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4798_ _0935_ _0941_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6468_ _2571_ _2574_ _2582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6304__A1 ci_adder.uut_simple_neuron.x3\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9256_ _0149_ net50 ci_adder.uut_simple_neuron.titan_id_6\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6399_ _2443_ _2511_ _2514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_9187_ _0220_ net76 ci_adder.uut_simple_neuron.titan_id_3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5419_ _1151_ _1559_ _1560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_8207_ ci_adder.output_val_internal\[31\] ci_adder.output_val_internal\[23\] ci_adder.output_val_internal\[15\]
+ ci_adder.output_val_internal\[7\] _3964_ _3961_ _4032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_100_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8138_ ci_adder.output_val_internal\[24\] ci_adder.output_val_internal\[16\] ci_adder.output_val_internal\[8\]
+ ci_adder.output_val_internal\[0\] _3964_ _3961_ _3970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8069_ internal_ih.byte5\[6\] internal_ih.byte4\[6\] _3919_ _3928_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8532__A2 _4235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9028__CLK net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8296__A1 _3645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6846__A2 ci_adder.uut_simple_neuron.x3\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9178__CLK net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4609__A1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8036__S _3908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5034__A1 ci_adder.uut_simple_neuron.x2\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8071__I1 internal_ih.byte4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5770_ _1895_ _1897_ _1898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_8_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4721_ _0877_ _0878_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_126_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4652_ _0766_ _0787_ ci_adder.uut_simple_neuron.x2\[8\] _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_72_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8523__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7440_ ci_adder.uut_simple_neuron.x0\[3\] _3452_ _3453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_126_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4583_ _0724_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7371_ _3397_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9110_ _0175_ net60 ci_adder.uut_simple_neuron.titan_id_0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6322_ _2398_ _2438_ _2439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8287__A1 _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6253_ _2049_ _2370_ _2371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9041_ ci_adder.input_memory\[1\]\[9\] net65 ci_adder.uut_simple_neuron.titan_id_1\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4848__A1 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5204_ _0717_ ci_adder.uut_simple_neuron.x2\[24\] _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6184_ _2300_ _2302_ _2303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout87_I net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5135_ _0870_ _1241_ _1283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5066_ _0831_ _1080_ _1214_ _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_84_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8695__CLK net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8173__C _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8825_ _0372_ net21 internal_ih.byte5\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5968_ _2047_ _2090_ _2091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5576__A2 ci_adder.uut_simple_neuron.x3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8756_ _0303_ net65 ci_adder.uut_simple_neuron.x2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_51_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4919_ _1070_ _1071_ _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7707_ _3502_ _3503_ _3670_ _3679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5899_ _2008_ _2010_ _2023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8687_ ci_adder.stream_o\[28\] ci_adder.output_memory\[28\] _4334_ _4343_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7638_ _1676_ _3617_ _3622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7569_ ci_adder.uut_simple_neuron.x0\[24\] ci_adder.uut_simple_neuron.x0\[25\] _3561_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_15_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9308_ _0569_ net45 ci_adder.stream_o\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9320__CLK net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8278__A1 _3608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9239_ _0103_ net84 ci_adder.uut_simple_neuron.titan_id_5\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8450__A1 _4165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6940_ _3038_ _3039_ _3040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5255__A1 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6871_ _2978_ _2979_ _2980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5822_ _1730_ _1948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8610_ _4257_ _4296_ _4298_ _4299_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5753_ _1878_ _1880_ _1881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_66_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8541_ _3524_ ci_adder.input_memory\[1\]\[17\] ci_adder.uut_simple_neuron.x2\[17\]
+ ci_adder.uut_simple_neuron.x3\[17\] _4206_ _4207_ _4243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_60_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4704_ _0860_ _0863_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_60_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5684_ _1768_ _1779_ _1814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8472_ ci_adder.output_val_internal\[4\] _4170_ _4187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4635_ _0797_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7423_ ci_adder.uut_simple_neuron.titan_id_1\[30\] ci_adder.uut_simple_neuron.titan_id_0\[30\]
+ _3441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4566_ _0724_ _0730_ _0731_ _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7354_ ci_adder.uut_simple_neuron.titan_id_1\[18\] ci_adder.uut_simple_neuron.titan_id_0\[18\]
+ _3383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6305_ _2250_ _2366_ _2421_ _2422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9024_ _0507_ net28 ci_adder.input_memory\[1\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7285_ _3311_ _3314_ _3324_ _3325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4497_ _0675_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6236_ _1999_ _2143_ _2354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7483__A2 ci_adder.uut_simple_neuron.x0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6167_ _0163_ _2285_ _2286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_90_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _1055_ _1264_ _1265_ _1266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8432__A1 internal_ih.spi_rx_byte_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6098_ _2023_ _2064_ _2115_ _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5246__A1 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5049_ _1138_ _1173_ _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5549__A2 _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8404__S _4139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8808_ _0355_ net23 internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8739_ _0286_ net42 internal_ih.spi_rx_byte_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8499__A1 _4165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8710__CLK net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5721__A2 _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6737__A1 _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8577__I2 ci_adder.uut_simple_neuron.x2\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4420_ _0602_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_112_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5472__I ci_adder.uut_simple_neuron.x2\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4351_ internal_ih.received_byte_count\[0\] _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_22_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7465__A2 _3470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7070_ _3146_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6021_ ci_adder.uut_simple_neuron.x3\[14\] _2099_ _2142_ _2143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__5476__A1 _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7217__A2 ci_adder.uut_simple_neuron.titan_id_5\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5228__A1 _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7972_ _3825_ _3877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6923_ ci_adder.uut_simple_neuron.titan_id_4\[7\] ci_adder.uut_simple_neuron.titan_id_3\[7\]
+ _3025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8017__I1 internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6854_ _2304_ _2901_ _2963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7776__I0 _3736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout38 net39 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout27 net40 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout16 net40 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_119_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5805_ _1867_ _1930_ _1931_ _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6785_ _2666_ _2894_ _2895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout49 net53 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5736_ _1831_ _1856_ _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8524_ _4211_ _4226_ _4228_ _4229_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5667_ _1772_ _1778_ _1797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8455_ ci_adder.uut_simple_neuron.x0\[1\] ci_adder.input_memory\[1\]\[1\] _0715_
+ _1676_ _4166_ _4167_ _4173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_79_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4618_ _0757_ _0777_ _0776_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7406_ ci_adder.uut_simple_neuron.titan_id_1\[27\] ci_adder.uut_simple_neuron.titan_id_0\[27\]
+ _3425_ _3426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5598_ ci_adder.uut_simple_neuron.x3\[5\] ci_adder.uut_simple_neuron.x3\[6\] _1731_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_8386_ _3667_ _4117_ _4130_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_92_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4549_ _0711_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7337_ _3369_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7268_ _3307_ _3309_ _3310_ _3311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_110_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6219_ _2335_ _2336_ _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9007_ _0490_ net58 ci_adder.input_memory\[1\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7208__A2 ci_adder.uut_simple_neuron.titan_id_5\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7199_ _3253_ _3254_ _3255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5219__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4690__A2 ci_adder.uut_simple_neuron.x2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6967__A1 ci_adder.uut_simple_neuron.titan_id_4\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_101_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8567__S1 _4253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8309__S _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4433__A2 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8044__S _3908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6570_ _2681_ _2682_ _2683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_4_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5521_ _1602_ _1652_ _1659_ _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_41_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8240_ _4050_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5452_ _1592_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7930__I0 _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5383_ _1340_ _1524_ _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4403_ internal_ih.byte4\[4\] _0623_ _0620_ internal_ih.byte0\[4\] _0626_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8171_ ci_adder.output_val_internal\[27\] ci_adder.output_val_internal\[19\] ci_adder.output_val_internal\[11\]
+ ci_adder.output_val_internal\[3\] _3964_ _3961_ _4000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_112_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7122_ ci_adder.uut_simple_neuron.titan_id_2\[8\] ci_adder.uut_simple_neuron.titan_id_5\[8\]
+ _3190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7053_ ci_adder.uut_simple_neuron.titan_id_4\[29\] ci_adder.uut_simple_neuron.titan_id_3\[29\]
+ _3133_ _3134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_74_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6004_ _1765_ _1769_ _2126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4546__I _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7610__A2 _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5621__A1 ci_adder.uut_simple_neuron.x3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7955_ _3868_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6906_ ci_adder.uut_simple_neuron.titan_id_4\[5\] ci_adder.uut_simple_neuron.titan_id_3\[5\]
+ _3011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7886_ internal_ih.received_byte_count\[2\] _3827_ _3829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6837_ _2944_ _2945_ _2946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_59_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6768_ _2842_ _2856_ _2877_ _2878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5924__A2 ci_adder.uut_simple_neuron.x3\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8507_ _4214_ _4215_ _4216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6699_ ci_adder.uut_simple_neuron.x3\[25\] _2735_ _2810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5719_ _1841_ _1847_ _1848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_115_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7677__A2 _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8438_ _3959_ _4157_ _3977_ _4158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8369_ _3625_ _4117_ _4121_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9061__CLK net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5860__A1 _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8779__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8485__S0 _4166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7968__S _3840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5612__A1 _1735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5915__A2 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7668__A2 _3645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8180__I3 ci_adder.output_val_internal\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4654__A2 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4366__I _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5603__A1 _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4952_ _1034_ _1068_ _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7740_ ci_adder.uut_simple_neuron.x0\[18\] _3695_ _3706_ _3599_ _3707_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4883_ _0965_ _0968_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7671_ _3608_ _3647_ _3648_ _3649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6622_ _2732_ _2733_ _2734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6553_ _2538_ _2665_ _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9084__CLK net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6484_ _2474_ _2538_ _2598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5504_ _1641_ _1642_ _1643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9272_ _0136_ net74 ci_adder.uut_simple_neuron.titan_id_6\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5435_ _1568_ _1575_ _1576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8223_ ci_adder.uut_simple_neuron.titan_id_6\[5\] _4042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5366_ _1421_ _1507_ _1508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8154_ _3960_ _3984_ _3985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5297_ _1401_ _1438_ _1439_ _1440_ _1441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_7105_ _3175_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8085_ _3936_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8921__CLK net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7036_ ci_adder.uut_simple_neuron.titan_id_4\[26\] ci_adder.uut_simple_neuron.titan_id_3\[26\]
+ _3118_ _3119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7788__S _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8987_ _0470_ net28 ci_adder.uut_simple_neuron.x0\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_78_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7938_ _3691_ _1011_ _3855_ _3860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_2_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5070__A2 _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8395__I0 _3691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8412__S _4139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7869_ _3805_ _3813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_21_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_76_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5570__I _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6086__A1 _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5833__A1 ci_adder.uut_simple_neuron.x3\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4636__A2 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_85_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8322__S _4091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6561__A2 _2673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_94_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8689__I1 ci_adder.output_memory\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5220_ _1329_ _1330_ _1365_ _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8944__CLK net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5151_ _1151_ _1276_ _1297_ _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6077__A1 _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5082_ _1089_ _1181_ _1230_ _1055_ _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_71_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8910_ _0038_ net12 ci_adder.value_i\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8449__S0 _4166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8841_ _0388_ net23 internal_ih.byte7\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8772_ _0319_ net71 ci_adder.uut_simple_neuron.x2\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5984_ _2103_ _2106_ _2107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7723_ _3691_ _2050_ _3692_ _3693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout32_I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4935_ _1081_ _1087_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6001__A1 _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4866_ _0970_ _0971_ _0969_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_82_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7654_ ci_adder.value_i\[4\] _3608_ _3635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6605_ _2715_ _2716_ _2717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6552__A2 ci_adder.uut_simple_neuron.x3\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4797_ _0927_ _0951_ _0952_ _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7585_ ci_adder.uut_simple_neuron.x0\[26\] ci_adder.uut_simple_neuron.x0\[27\] _3574_
+ _3575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_6_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6536_ _2588_ _2627_ _2649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4563__A1 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8031__I _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6467_ _2579_ _2580_ _2581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6304__A2 _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9255_ _0138_ net50 ci_adder.uut_simple_neuron.titan_id_6\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6398_ _2510_ _2507_ _2511_ _2446_ _2512_ _2513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_113_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9186_ _0219_ net77 ci_adder.uut_simple_neuron.titan_id_3\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5418_ _1084_ _1558_ _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8206_ _3963_ ci_adder.stream_o\[7\] ci_adder.stream_o\[23\] _3965_ _4030_ _4031_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5349_ _1477_ _1491_ _1492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8137_ _3963_ ci_adder.stream_o\[0\] ci_adder.stream_o\[16\] _3965_ _3968_ _3969_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__6068__A1 _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8068_ _3927_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7019_ ci_adder.uut_simple_neuron.titan_id_4\[24\] ci_adder.uut_simple_neuron.titan_id_3\[24\]
+ _3105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8817__CLK net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8612__S0 _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8296__A2 _4071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6059__A1 _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4720_ _0877_ _0878_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4651_ ci_adder.uut_simple_neuron.x2\[6\] _0809_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7731__A1 _3524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4582_ _0714_ _0741_ _0742_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7370_ _3395_ _3396_ _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_52_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6321_ _2400_ _2437_ _2438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8531__I0 ci_adder.uut_simple_neuron.x0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8287__A2 _4071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6252_ _2051_ _2199_ _2370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9040_ ci_adder.input_memory\[1\]\[8\] net65 ci_adder.uut_simple_neuron.titan_id_1\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9122__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6183_ _2200_ _2301_ _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5203_ _0711_ _1348_ _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5134_ _1213_ _1240_ _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9272__CLK net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5065_ _0831_ _0939_ _1082_ _1214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_84_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8824_ _0371_ net21 internal_ih.byte5\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5967_ _1919_ _2052_ _2090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8755_ _0302_ net65 ci_adder.uut_simple_neuron.x2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_51_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4918_ _0993_ _1063_ _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4784__A1 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7706_ _3678_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8686_ _4342_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5898_ _2014_ _2022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_47_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7637_ _0065_ _3619_ _3620_ _3621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__6525__A2 _2638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4849_ _0874_ _0909_ _0931_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_7568_ _3560_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6519_ _1726_ _1728_ _2633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7499_ ci_adder.uut_simple_neuron.x0\[12\] _3502_ _3503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9307_ _0568_ net46 ci_adder.stream_o\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9238_ _0102_ net84 ci_adder.uut_simple_neuron.titan_id_5\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9169_ _0202_ net87 ci_adder.uut_simple_neuron.titan_id_3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9145__CLK net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6870_ _1882_ _2912_ _2979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5821_ _1913_ _1925_ _1946_ _1947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7952__A1 ci_adder.uut_simple_neuron.x2\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ ci_adder.uut_simple_neuron.x3\[9\] _1879_ _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_22_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8540_ ci_adder.output_memory\[17\] _4212_ _4242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4703_ _0830_ _0861_ _0862_ _0841_ _0804_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_17_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5683_ _1795_ _1799_ _1812_ _1813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8471_ _4165_ _4185_ _4186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4634_ _0782_ _0783_ _0796_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_71_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7422_ _3415_ _3423_ _3435_ _3439_ _3440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_32_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4565_ _0724_ ci_adder.uut_simple_neuron.x2\[4\] _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7353_ _3382_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6304_ ci_adder.uut_simple_neuron.x3\[20\] _2365_ _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_69_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4549__I _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9023_ _0506_ net28 ci_adder.input_memory\[1\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7284_ ci_adder.uut_simple_neuron.titan_id_1\[5\] ci_adder.uut_simple_neuron.titan_id_0\[5\]
+ _3324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4496_ internal_ih.byte3\[0\] _0670_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_31_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6235_ _2294_ _2310_ _2352_ _2353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6166_ _1871_ _1886_ _2285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6097_ _2215_ _2217_ _2218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_90_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _1224_ _1228_ _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5048_ _1194_ _1197_ _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__9018__CLK net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8196__A1 _3966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8807_ _0354_ net23 internal_ih.byte3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_40_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6999_ _3088_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6746__A2 _2856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9168__CLK net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8738_ _0285_ net43 internal_ih.spi_rx_byte_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_47_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8669_ _4333_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8499__A2 _4208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8420__S _4139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6682__A1 _2720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8187__A1 _3966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8577__I3 _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4748__A1 ci_adder.uut_simple_neuron.x2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8330__S _4091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5173__A1 _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4350_ internal_ih.received_byte_count\[4\] internal_ih.received_byte_count\[7\]
+ internal_ih.received_byte_count\[6\] _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_39_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6673__A1 _2720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6020_ _2050_ _2098_ _2142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5476__A2 ci_adder.uut_simple_neuron.x2\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6425__A1 _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7971_ _3876_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6922_ _3024_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8178__A1 _3966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6853_ ci_adder.uut_simple_neuron.x3\[30\] _2356_ _2961_ _2962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_89_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9310__CLK net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5804_ _1869_ _1890_ _1931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7776__I1 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout28 net31 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_9_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout17 net18 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6784_ _2892_ _2893_ _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout39 net40 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5735_ _1824_ _1861_ _1862_ _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_91_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout9_I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8523_ ci_adder.output_val_internal\[13\] _4203_ _4229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5666_ _1770_ _1796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8454_ ci_adder.output_memory\[1\] _4163_ _4172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_79_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4617_ _0780_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7405_ _3419_ _3424_ _3425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5597_ ci_adder.uut_simple_neuron.x3\[3\] _1712_ _1729_ _1730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_8385_ ci_adder.input_memory\[1\]\[10\] _4118_ _4130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4548_ _0716_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7336_ _3366_ _3368_ _3369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4479_ internal_ih.byte2\[0\] _0659_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7267_ ci_adder.uut_simple_neuron.titan_id_1\[4\] ci_adder.uut_simple_neuron.titan_id_0\[4\]
+ _3310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6218_ _2281_ _2287_ _2336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9006_ _0489_ net59 ci_adder.input_memory\[1\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7198_ ci_adder.uut_simple_neuron.titan_id_2\[22\] ci_adder.uut_simple_neuron.titan_id_5\[22\]
+ _3254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6149_ _2172_ _2214_ _2269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8169__A1 _3966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7916__A1 _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4902__A1 _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6655__A1 _2694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_19_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4969__A1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7907__A1 _3616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5520_ _1487_ _1658_ _1659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5451_ _1588_ _1591_ _1592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_41_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5382_ _1263_ _1523_ _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4402_ _0625_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8170_ _3963_ ci_adder.stream_o\[3\] ci_adder.stream_o\[19\] _3965_ _3998_ _3999_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_112_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7121_ _3189_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7052_ _3110_ _3111_ _3127_ _3132_ _3133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__6646__A1 _2147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6003_ _2123_ _2124_ _2125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_105_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout62_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7954_ _3733_ ci_adder.uut_simple_neuron.x2\[23\] _3840_ _3868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5621__A2 ci_adder.uut_simple_neuron.x3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6905_ _3006_ _3008_ _3009_ _3010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_82_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7885_ internal_ih.received_byte_count\[2\] _3827_ _3828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6836_ _2876_ _2935_ _2945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_114_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6767_ _2801_ _2841_ _2877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_57_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8850__CLK net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5718_ _1754_ _1846_ _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_73_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8506_ ci_adder.uut_simple_neuron.x0\[10\] ci_adder.input_memory\[1\]\[10\] ci_adder.uut_simple_neuron.x2\[10\]
+ ci_adder.uut_simple_neuron.x3\[10\] _4206_ _4207_ _4215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_17_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6698_ ci_adder.uut_simple_neuron.x3\[26\] ci_adder.uut_simple_neuron.x3\[27\] _2809_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5649_ _1768_ _1779_ _1780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8437_ internal_ih.spi_rx_byte_i\[1\] _3812_ _3966_ _4157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8368_ ci_adder.input_memory\[1\]\[2\] _4118_ _4121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7319_ ci_adder.uut_simple_neuron.titan_id_1\[12\] ci_adder.uut_simple_neuron.titan_id_0\[12\]
+ _3355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_123_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8299_ _3479_ _4072_ _4082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8485__S1 _4167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5128__A1 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6876__A1 _2921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5300__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8723__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8055__S _3919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7979__I1 internal_ih.spi_rx_byte_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5603__A2 _1715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8873__CLK net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4951_ _1064_ _1067_ _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4882_ _1000_ _1023_ _1035_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7670_ _3469_ _3638_ _3470_ _3648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6621_ _2538_ _2665_ _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9229__CLK net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6552_ ci_adder.uut_simple_neuron.x3\[25\] ci_adder.uut_simple_neuron.x3\[26\] _2665_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8305__A1 _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6483_ _2474_ _2538_ _2597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5503_ _1602_ _1633_ _1642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9271_ _0135_ net81 ci_adder.uut_simple_neuron.titan_id_6\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5434_ _1573_ _1574_ _1575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8222_ _4041_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8153_ ci_adder.output_val_internal\[25\] ci_adder.output_val_internal\[17\] ci_adder.output_val_internal\[9\]
+ ci_adder.output_val_internal\[1\] _3964_ _3961_ _3984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_100_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5365_ _1463_ _1503_ _1507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7104_ _3173_ _3174_ _3175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_22_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8608__A2 _4297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5296_ _1400_ _1407_ _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8084_ internal_ih.byte6\[5\] internal_ih.byte5\[5\] _3930_ _3936_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7035_ _3110_ _3111_ _3117_ _3114_ _3118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7868__I _3811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8986_ _0469_ net25 ci_adder.uut_simple_neuron.x0\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_78_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7937_ _3859_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7868_ _3811_ _3812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6819_ _1871_ _2928_ _2929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8544__A1 _4211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7799_ ci_adder.value_i\[28\] _3659_ _3756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8746__CLK net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5833__A2 ci_adder.uut_simple_neuron.x3\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8896__CLK net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5597__A1 ci_adder.uut_simple_neuron.x3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8535__A1 ci_adder.output_memory\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5150_ _1110_ _1275_ _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6077__A2 ci_adder.uut_simple_neuron.x3\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5081_ _1124_ _1162_ _1230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_71_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8449__S1 _4167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8840_ _0387_ net21 internal_ih.byte7\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5983_ _2105_ _2106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8771_ _0318_ net73 ci_adder.uut_simple_neuron.x2\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9051__CLK net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4934_ _1084_ _1086_ _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7722_ _3611_ _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_59_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_82_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4865_ _0970_ _0969_ _0971_ _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_fanout25_I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7653_ _3452_ _3627_ _3634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6604_ _2706_ _2711_ _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4796_ _0930_ _0943_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_74_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7584_ _3572_ _3573_ _3574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6535_ _2629_ _2637_ _2647_ _2648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9254_ _0127_ net51 ci_adder.uut_simple_neuron.titan_id_6\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6466_ _2517_ _2577_ _2580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8205_ _3966_ _4029_ _4030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6397_ _2389_ _2441_ _2504_ _2512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_9185_ _0218_ net76 ci_adder.uut_simple_neuron.titan_id_3\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5417_ _1263_ _1523_ _1557_ _1558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5512__A1 _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5348_ _1482_ _1490_ _1491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8136_ _3966_ _3967_ _3968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6068__A2 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8301__I1 ci_adder.uut_simple_neuron.x0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8067_ internal_ih.byte5\[5\] internal_ih.byte4\[5\] _3919_ _3927_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7018_ _3102_ _3103_ _3104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5279_ _1421_ _1423_ _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5579__A1 ci_adder.uut_simple_neuron.x3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8969_ _0452_ net56 ci_adder.uut_simple_neuron.x0\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8612__S1 _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5751__A1 ci_adder.uut_simple_neuron.x3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9074__CLK net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5756__I _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4650_ _0766_ _0787_ _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_44_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8911__CLK net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6320_ _2410_ _2436_ _2437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4581_ _0740_ _0732_ _0745_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6251_ _2245_ _2368_ _2369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6182_ _2250_ ci_adder.uut_simple_neuron.x3\[20\] _2301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_5202_ ci_adder.uut_simple_neuron.x2\[24\] _1348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_5133_ _0870_ _1280_ _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5064_ _1212_ _1190_ _1191_ _1156_ _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_84_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8823_ _0370_ net21 internal_ih.byte5\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4481__A1 internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _1750_ _2088_ _2089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8754_ _0301_ net82 ci_adder.uut_simple_neuron.x2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5981__A1 _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ _2021_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4917_ _1036_ _1062_ _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7705_ _3677_ ci_adder.uut_simple_neuron.x3\[12\] _3632_ _3678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8685_ ci_adder.stream_o\[27\] ci_adder.output_memory\[27\] _4334_ _4342_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4848_ _0831_ _1001_ _1002_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_62_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7636_ ci_adder.value_i\[1\] _3599_ _3620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_105_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4779_ ci_adder.uut_simple_neuron.x2\[6\] _0809_ _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7567_ _3556_ _3559_ _3560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7881__I _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9306_ _0567_ net47 ci_adder.stream_o\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6518_ _2630_ _2631_ _2632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_95_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7498_ ci_adder.uut_simple_neuron.x0\[13\] _3502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_43_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ _2040_ _2056_ _2564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6289__A2 _2356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9237_ _0101_ net83 ci_adder.uut_simple_neuron.titan_id_5\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9168_ _0201_ net87 ci_adder.uut_simple_neuron.titan_id_3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8119_ internal_ih.current_instruction\[6\] _3947_ _3954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__9097__CLK net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8418__S _4139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9099_ _0194_ net62 ci_adder.uut_simple_neuron.titan_id_0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5972__A1 ci_adder.uut_simple_neuron.x3\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7961__A2 _3841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8597__S0 _4252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7713__A2 _3659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8521__S0 _4206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8127__I _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5820_ _1911_ _1926_ _1946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8063__S _3919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5751_ ci_adder.uut_simple_neuron.x3\[10\] ci_adder.uut_simple_neuron.x3\[11\] _1879_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__7952__A2 _3846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _0832_ _0839_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_60_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8470_ _3452_ ci_adder.input_memory\[1\]\[4\] ci_adder.uut_simple_neuron.x2\[4\]
+ ci_adder.uut_simple_neuron.x3\[4\] _4166_ _4167_ _4185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_8_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5682_ _1808_ _1811_ _1812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_60_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7421_ _3438_ _3439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5715__A1 ci_adder.uut_simple_neuron.x3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4633_ _0786_ _0795_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4564_ _0722_ ci_adder.uut_simple_neuron.x2\[4\] _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7352_ _3380_ _3381_ _3382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_52_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6303_ _2245_ _2368_ _2419_ _2420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7283_ _3323_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7468__A1 _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout92_I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6234_ _2296_ _2309_ _2352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9022_ _0505_ net28 ci_adder.input_memory\[1\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4495_ _0674_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8807__CLK net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6165_ _2282_ _2283_ _2284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6096_ _2162_ _2160_ _2216_ _2217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_90_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _1224_ _1228_ _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5047_ _0996_ _1195_ _1196_ _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8957__CLK net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7640__A1 ci_adder.uut_simple_neuron.x0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4454__A1 internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6998_ ci_adder.uut_simple_neuron.titan_id_4\[20\] ci_adder.uut_simple_neuron.titan_id_3\[20\]
+ _3087_ _3088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_95_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8806_ _0353_ net40 internal_ih.byte2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5949_ _2017_ _2020_ _2067_ _2069_ _2072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_94_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8737_ _0284_ net43 internal_ih.spi_rx_byte_i\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8668_ ci_adder.stream_o\[19\] ci_adder.output_memory\[19\] _4323_ _4333_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7619_ _0700_ _3597_ _3604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8599_ ci_adder.output_val_internal\[27\] _4249_ _4291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6131__A1 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6434__A2 _2364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7631__A1 ci_adder.value_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9112__CLK net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7698__A1 _3629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_117_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8498__I0 ci_adder.uut_simple_neuron.x0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8111__A2 _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6122__A1 _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7970_ _3768_ ci_adder.uut_simple_neuron.x2\[31\] _3840_ _3876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6921_ _3022_ _3023_ _3024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6852_ _1695_ _2952_ _2960_ _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8422__I0 _3757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5803_ _1869_ _1890_ _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout29 net31 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout18 net40 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_119_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6783_ ci_adder.uut_simple_neuron.x3\[29\] _2812_ _2893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8522_ _4214_ _4227_ _4228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5734_ _1859_ _1860_ _1857_ _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_45_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5665_ _1793_ _1794_ _1795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8453_ _4162_ _4164_ _4169_ _4171_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_79_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4616_ _0761_ _0779_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8384_ _4129_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7404_ ci_adder.uut_simple_neuron.titan_id_1\[27\] ci_adder.uut_simple_neuron.titan_id_0\[27\]
+ _3424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5596_ ci_adder.uut_simple_neuron.x3\[4\] ci_adder.uut_simple_neuron.x3\[5\] _1729_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7335_ _3367_ _3368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4547_ _0710_ _0715_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6113__A1 _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4478_ _0665_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7266_ ci_adder.uut_simple_neuron.titan_id_1\[4\] ci_adder.uut_simple_neuron.titan_id_0\[4\]
+ _3309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6217_ _2284_ _2286_ _2335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7197_ _3243_ _3248_ _3249_ _3251_ _3252_ _3253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_9005_ _0488_ net59 ci_adder.input_memory\[1\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7861__A1 internal_ih.spi_rx_byte_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6148_ _2265_ _2267_ _2268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__9135__CLK net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6079_ ci_adder.uut_simple_neuron.x3\[18\] _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4427__B2 internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7916__A2 _3841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5927__A1 ci_adder.uut_simple_neuron.x3\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6352__A1 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__A2 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7852__A1 _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4666__A1 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4418__B2 internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4969__A2 _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8404__I0 _3713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7907__A2 _3841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5450_ _1589_ _1590_ _1591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9008__CLK net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4401_ internal_ih.byte4\[3\] _0623_ _0620_ internal_ih.byte0\[3\] _0625_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5381_ _1480_ _1481_ _1522_ _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_1_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7120_ _3187_ _3188_ _3189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_120_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7051_ ci_adder.uut_simple_neuron.titan_id_4\[28\] ci_adder.uut_simple_neuron.titan_id_3\[28\]
+ _3126_ _3129_ _3131_ _3132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6646__A2 _2673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7843__A1 _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6002_ _1750_ _2088_ _2124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_74_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4409__A1 internal_ih.byte4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4409__B2 internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7953_ _3728_ _3842_ _3867_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout55_I net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5082__B2 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6904_ ci_adder.uut_simple_neuron.titan_id_4\[4\] ci_adder.uut_simple_neuron.titan_id_3\[4\]
+ _3009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7884_ _3823_ _3826_ _3827_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6835_ _2879_ _2934_ _2944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6582__A1 _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6766_ _2844_ _2855_ _2875_ _2876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_92_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5717_ _1843_ _1845_ _1846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_18_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8505_ _0704_ _4214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_115_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6697_ _2540_ _2737_ _2807_ _2808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5648_ _1770_ _1772_ _1778_ _1779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8436_ _4156_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5579_ ci_adder.uut_simple_neuron.x3\[3\] _1712_ _1713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_4
XFILLER_0_20_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8367_ _3621_ _4117_ _4120_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7318_ _3350_ _3351_ _3352_ _3353_ _3354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_8298_ _3650_ _4071_ _4081_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7249_ ci_adder.uut_simple_neuron.titan_id_2\[30\] ci_adder.uut_simple_neuron.titan_id_5\[30\]
+ _3297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_99_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8426__S _4116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5073__A1 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5128__A2 _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9300__CLK net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8336__S _4091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4950_ _1072_ _1102_ _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4811__A1 _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4881_ _1019_ _1022_ _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6620_ ci_adder.uut_simple_neuron.x3\[25\] ci_adder.uut_simple_neuron.x3\[26\] _2732_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8071__S _3919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6551_ _2474_ _2600_ _2663_ _2664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_61_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5502_ _1629_ _1632_ _1641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8305__A2 _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6316__A1 _1962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6482_ _2367_ _2594_ _2595_ _2596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5119__A2 ci_adder.uut_simple_neuron.x2\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9270_ _0134_ net81 ci_adder.uut_simple_neuron.titan_id_6\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5433_ ci_adder.uut_simple_neuron.x2\[29\] _1532_ _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8221_ ci_adder.uut_simple_neuron.titan_id_6\[4\] _4041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5364_ _1506_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8152_ _3963_ ci_adder.stream_o\[1\] ci_adder.stream_o\[17\] _3965_ _3982_ _3983_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__4838__I _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7103_ ci_adder.uut_simple_neuron.titan_id_2\[7\] ci_adder.uut_simple_neuron.titan_id_5\[7\]
+ _3174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5295_ _1402_ _1405_ _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8083_ _3935_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7034_ ci_adder.uut_simple_neuron.titan_id_4\[26\] ci_adder.uut_simple_neuron.titan_id_3\[26\]
+ _3117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8985_ _0468_ net26 ci_adder.uut_simple_neuron.x0\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_7936_ _3685_ ci_adder.uut_simple_neuron.x2\[14\] _3855_ _3859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_65_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7867_ _3807_ _3810_ internal_ih.instruction_received _3811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_38_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _1876_ _1886_ _2928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7798_ ci_adder.uut_simple_neuron.x0\[28\] _3753_ _3614_ _3755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6749_ _2723_ _2860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_107_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6307__A1 ci_adder.uut_simple_neuron.x3\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8419_ _4147_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8535__A2 _4212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8299__A1 _3479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5080_ _1016_ _1224_ _1228_ _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_71_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8840__CLK net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8471__A1 _4165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5285__A1 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4393__I _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5982_ _1843_ _2104_ _2105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8770_ _0317_ net73 ci_adder.uut_simple_neuron.x2\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_63_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8990__CLK net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4933_ _1055_ _1085_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7721_ _3619_ _3688_ _3689_ _3690_ _3691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_82_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4864_ _1003_ _1010_ _1018_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_74_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7652_ _3633_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6603_ _2713_ _2714_ _2640_ _2705_ _2715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_105_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4795_ _0930_ _0943_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_62_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7583_ _3569_ _3570_ _3573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout18_I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6534_ _2632_ _2636_ _2647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6465_ _2518_ _2575_ _2579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9253_ _0119_ net71 ci_adder.uut_simple_neuron.titan_id_5\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5416_ _1340_ _1524_ _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8204_ _3962_ ci_adder.stream_o\[15\] _4029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6396_ _2442_ _2504_ _2511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_113_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9184_ _0217_ net77 ci_adder.uut_simple_neuron.titan_id_3\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5512__A2 ci_adder.uut_simple_neuron.x2\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5347_ _1483_ _1489_ _1490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8135_ _3962_ ci_adder.stream_o\[8\] _3967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5278_ _1367_ _1422_ _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8066_ _3926_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7017_ _3099_ _3100_ _3103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8065__I1 internal_ih.byte4\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8968_ _0451_ net58 ci_adder.uut_simple_neuron.x0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7919_ _0766_ _3842_ _3850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8899_ _0058_ net12 ci_adder.value_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8503__I _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5751__A2 ci_adder.uut_simple_neuron.x3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8863__CLK net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8205__A1 _3966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_122_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8508__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4580_ _0724_ _0722_ ci_adder.uut_simple_neuron.x2\[4\] _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_65_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6250_ _2364_ _2367_ _2368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8531__I2 _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6181_ ci_adder.uut_simple_neuron.x3\[17\] _2251_ _2299_ _2300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5201_ _0713_ _1316_ _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5132_ _1249_ _1279_ _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5258__A1 ci_adder.uut_simple_neuron.x2\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5063_ _1180_ _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8822_ _0369_ net16 internal_ih.byte4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4481__A2 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5965_ _1756_ _2087_ _2088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8753_ _0300_ net86 ci_adder.uut_simple_neuron.x2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_51_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5896_ _2017_ _2020_ _2021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5981__A2 _1958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4916_ _1069_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7704_ _3674_ _3676_ _3677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8684_ _4341_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4847_ _0965_ _0968_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_28_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7635_ _3608_ _3619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_117_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4778_ _0766_ _0787_ ci_adder.uut_simple_neuron.x2\[8\] _0909_ _0935_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7566_ _3553_ _3557_ _3558_ _3552_ _3559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_9305_ _0566_ net46 ci_adder.stream_o\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6517_ _2560_ _2566_ _2631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7497_ _3501_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6448_ _2561_ _2486_ _2562_ _2563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_95_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9236_ _0100_ net88 ci_adder.uut_simple_neuron.titan_id_5\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6379_ _1989_ _2004_ _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9167_ _0227_ net87 ci_adder.uut_simple_neuron.titan_id_3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8118_ _3953_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9098_ _0193_ net61 ci_adder.uut_simple_neuron.titan_id_0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6997__A1 _3083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8049_ _3917_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8038__I1 internal_ih.byte2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_104_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5972__A2 _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8597__S1 _4253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7740__C _3599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8521__S1 _4207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9191__CLK net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8029__I1 internal_ih.byte2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8344__S _4070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7788__I0 _3746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5963__A2 _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5750_ ci_adder.uut_simple_neuron.x3\[8\] _1844_ _1877_ _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5681_ _1810_ _1811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4701_ _0832_ _0839_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4632_ _0773_ _0794_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7420_ _3430_ _3436_ _3435_ _3426_ _3437_ _3438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5715__A2 ci_adder.uut_simple_neuron.x3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4563_ _0718_ _0720_ _0728_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_69_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7351_ ci_adder.uut_simple_neuron.titan_id_1\[18\] ci_adder.uut_simple_neuron.titan_id_0\[18\]
+ _3381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6302_ _2364_ _2418_ _2419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7282_ _3321_ _3322_ _3323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7468__A2 _3470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4494_ internal_ih.byte2\[7\] _0670_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6233_ _2344_ _2350_ _2351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9021_ _0504_ net29 ci_adder.input_memory\[1\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6164_ _1841_ _2241_ _2283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout85_I net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6095_ _2156_ _2159_ _2216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _1260_ _1262_ _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5046_ _1149_ _1170_ _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6997_ _3083_ _3085_ _3086_ _3087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_79_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8805_ _0352_ net17 internal_ih.byte2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5948_ _2071_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8736_ _0283_ net43 internal_ih.spi_rx_byte_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_47_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5879_ _1774_ _2003_ _2004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8667_ _4332_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7618_ _3599_ _3601_ _3602_ _3603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_8598_ _4260_ _4289_ _4290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7549_ ci_adder.uut_simple_neuron.x0\[19\] _3539_ _3544_ _3545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9064__CLK net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4390__B2 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9219_ _0085_ net30 ci_adder.uut_simple_neuron.titan_id_2\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6131__A2 _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8901__CLK net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7631__A2 _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5642__A1 ci_adder.uut_simple_neuron.x3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7942__I0 _3703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8498__I1 ci_adder.input_memory\[1\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4381__B2 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7870__A2 internal_ih.spi_rx_byte_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6920_ ci_adder.uut_simple_neuron.titan_id_4\[7\] ci_adder.uut_simple_neuron.titan_id_3\[7\]
+ _3023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8074__S _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6851_ _2541_ _2956_ _2959_ _2960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_77_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5802_ _1904_ _1928_ _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_9_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout19 net21 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_119_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6782_ _2890_ _2891_ _2892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8521_ _3502_ ci_adder.input_memory\[1\]\[13\] ci_adder.uut_simple_neuron.x2\[13\]
+ ci_adder.uut_simple_neuron.x3\[13\] _4206_ _4207_ _4227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_57_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5733_ _1859_ _1860_ _1857_ _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9087__CLK net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5664_ _1681_ _1711_ _1675_ _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8452_ ci_adder.output_val_internal\[0\] _4170_ _4171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5595_ _1681_ _1714_ _1727_ _1728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_4615_ _0776_ _0778_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_79_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8383_ _3661_ ci_adder.input_memory\[1\]\[9\] _4122_ _4129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7403_ _3416_ _3421_ _3423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4546_ _0714_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7334_ ci_adder.uut_simple_neuron.titan_id_1\[15\] ci_adder.uut_simple_neuron.titan_id_0\[15\]
+ _3367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4372__B2 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4477_ internal_ih.byte1\[7\] _0659_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8924__CLK net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7265_ _3308_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6216_ _2334_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7196_ ci_adder.uut_simple_neuron.titan_id_2\[21\] ci_adder.uut_simple_neuron.titan_id_5\[21\]
+ _3252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9004_ _0487_ net59 ci_adder.input_memory\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6147_ _2176_ _2213_ _2266_ _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_110_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5872__A1 ci_adder.uut_simple_neuron.x3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5624__A1 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6078_ _2050_ _2144_ _2198_ _2199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__4427__A2 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5029_ _1158_ _1166_ _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5927__A2 ci_adder.uut_simple_neuron.x3\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8719_ _0274_ net71 ci_adder.uut_simple_neuron.x3\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6352__A2 _2423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4363__A1 internal_ih.current_instruction\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5863__A1 _1754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4418__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8652__I1 ci_adder.output_memory\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_19_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8947__CLK net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4400_ _0624_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5380_ _1447_ _1479_ _1522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_50_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8069__S _3919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8340__I0 _3757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7050_ _3130_ _3131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6001_ _1756_ _2087_ _2123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4409__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8643__I1 ci_adder.output_memory\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7952_ ci_adder.uut_simple_neuron.x2\[22\] _3846_ _3867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_19_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6903_ ci_adder.uut_simple_neuron.titan_id_4\[4\] ci_adder.uut_simple_neuron.titan_id_3\[4\]
+ _3008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout48_I net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7883_ internal_ih.received_byte_count\[1\] _3822_ _3827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_119_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6834_ _2545_ _2941_ _2942_ _2943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6765_ _2847_ _2854_ _2875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5716_ ci_adder.uut_simple_neuron.x3\[8\] _1844_ _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_18_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8504_ ci_adder.output_memory\[10\] _4212_ _4213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6696_ _2734_ _2736_ _2807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8435_ _4154_ _4155_ _4156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_17_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5647_ _1713_ _1777_ _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_60_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7531__A1 ci_adder.uut_simple_neuron.x0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5578_ ci_adder.uut_simple_neuron.x3\[4\] ci_adder.uut_simple_neuron.x3\[5\] _1712_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_14_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8366_ ci_adder.input_memory\[1\]\[1\] _4118_ _4120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7317_ ci_adder.uut_simple_neuron.titan_id_1\[11\] ci_adder.uut_simple_neuron.titan_id_0\[11\]
+ _3353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8297_ _3470_ _4072_ _4081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4529_ _0697_ _0698_ ci_adder.address_i\[2\] _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7248_ _3292_ _3294_ _3295_ _3296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__9102__CLK net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5845__A1 _1945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4648__A2 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7179_ _3237_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_37_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A1 _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_46_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8241__I ci_adder.uut_simple_neuron.titan_id_6\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8322__I0 _3713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5836__A1 _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8389__I0 _3677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6013__A1 _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4880_ _1028_ _1031_ _1033_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_86_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_64_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6550_ _2538_ ci_adder.uut_simple_neuron.x3\[25\] _2663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_39_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5501_ _1640_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6481_ _2537_ _2540_ _2595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_76_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5432_ _1569_ _1570_ _1572_ _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_2_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8220_ _4040_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9125__CLK net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5363_ _1503_ _1505_ _1506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8151_ _3966_ _3981_ _3982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8313__I0 _3691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7102_ ci_adder.uut_simple_neuron.titan_id_2\[6\] ci_adder.uut_simple_neuron.titan_id_5\[6\]
+ _3172_ _3173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5827__A1 _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5294_ _1402_ _1405_ _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8082_ internal_ih.byte6\[4\] internal_ih.byte5\[4\] _3930_ _3935_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7033_ _3116_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6252__A1 _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8984_ _0467_ net26 ci_adder.uut_simple_neuron.x0\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7230__I _3280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7935_ _3858_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7866_ _3808_ _3809_ _3810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6817_ _2925_ _2926_ _2927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4566__A1 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7797_ ci_adder.uut_simple_neuron.x0\[28\] _3753_ _3754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6748_ _2797_ _2858_ _2859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6679_ _2710_ _2788_ _2790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6307__A2 _2423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8418_ _3746_ ci_adder.input_memory\[1\]\[26\] _4139_ _4147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8349_ _3963_ _3974_ _3975_ _4107_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5818__A1 _1682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9148__CLK net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8299__A2 _4072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9298__CLK net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5981_ _1845_ _1958_ _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_87_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4932_ _1011_ ci_adder.uut_simple_neuron.x2\[16\] _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8082__S _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7720_ ci_adder.value_i\[15\] _3659_ _3690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7651_ _3631_ ci_adder.uut_simple_neuron.x3\[3\] _3632_ _3633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6602_ _2520_ _2570_ _2714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6537__A2 _2638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4863_ _0978_ _1017_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4794_ _0922_ _0946_ _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7582_ ci_adder.uut_simple_neuron.x0\[25\] ci_adder.uut_simple_neuron.x0\[26\] _3572_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6533_ _2640_ _2642_ _2646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9321_ _0582_ net45 ci_adder.stream_o\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6464_ _2578_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9252_ _0117_ net71 ci_adder.uut_simple_neuron.titan_id_5\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5415_ _1554_ _1555_ _1556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8203_ _3979_ _4027_ _4028_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6395_ _2389_ _2441_ _2504_ _2510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_9183_ _0216_ net77 ci_adder.uut_simple_neuron.titan_id_3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5346_ _1487_ _1488_ _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8134_ _3964_ _3966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5277_ _1374_ _1376_ _1382_ _1369_ _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_8065_ internal_ih.byte5\[4\] internal_ih.byte4\[4\] _3919_ _3926_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8462__A2 _4170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7016_ ci_adder.uut_simple_neuron.titan_id_4\[23\] ci_adder.uut_simple_neuron.titan_id_3\[23\]
+ _3102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6225__A1 _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8967_ _0450_ net62 ci_adder.uut_simple_neuron.x0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_26_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7918_ _3641_ _3841_ _3849_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_54_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8898_ _0055_ net13 ci_adder.value_i\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7849_ _3770_ _3795_ _3796_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4778__A1 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7192__A2 ci_adder.uut_simple_neuron.titan_id_5\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8531__I3 _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6180_ _2200_ _2250_ _2299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5200_ _1314_ _1317_ _1345_ _1316_ _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_5131_ _1251_ _1256_ _1278_ _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5062_ _0993_ _1193_ _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5258__A2 ci_adder.uut_simple_neuron.x2\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8821_ _0368_ net16 internal_ih.byte4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9313__CLK net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4769__A1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8752_ _0299_ net73 ci_adder.uut_simple_neuron.x2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5964_ _1803_ _2055_ _2086_ _2087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_fanout30_I net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7703_ _3497_ _3663_ _3675_ _3614_ _3676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_118_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5895_ _1941_ _2018_ _2019_ _2020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_4915_ _1034_ _1068_ _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_51_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8683_ ci_adder.stream_o\[26\] ci_adder.output_memory\[26\] _4334_ _4341_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4846_ _0965_ _0968_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7634_ _3612_ _3616_ _3618_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7183__A2 ci_adder.uut_simple_neuron.titan_id_5\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7565_ ci_adder.uut_simple_neuron.x0\[22\] ci_adder.uut_simple_neuron.x0\[23\] _3558_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6516_ _2563_ _2565_ _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4777_ ci_adder.uut_simple_neuron.x2\[13\] _0932_ _0933_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9304_ _0565_ net46 ci_adder.stream_o\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7496_ _3497_ _3500_ _3501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6447_ _2043_ _2485_ _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_95_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9235_ _0099_ net85 ci_adder.uut_simple_neuron.titan_id_5\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6378_ _2492_ _2493_ _2494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9166_ _0226_ net87 ci_adder.uut_simple_neuron.titan_id_3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5329_ _1437_ _1455_ _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8117_ internal_ih.current_instruction\[5\] _3947_ _3953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_9097_ _0190_ net61 ci_adder.uut_simple_neuron.titan_id_0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8048_ internal_ih.byte4\[4\] internal_ih.byte3\[4\] _3908_ _3917_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8199__A1 _3811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8830__CLK net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4932__A1 _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4999__A1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7788__I1 ci_adder.uut_simple_neuron.x3\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5680_ _1690_ _1809_ _1810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4700_ _0845_ _0859_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_84_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4631_ _0792_ _0793_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4562_ _0709_ ci_adder.uut_simple_neuron.x2\[2\] _0722_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7350_ _3375_ _3377_ _3379_ _3380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_52_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ _2250_ _2366_ _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7281_ ci_adder.uut_simple_neuron.titan_id_1\[7\] ci_adder.uut_simple_neuron.titan_id_0\[7\]
+ _3322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4493_ _0673_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6232_ _2347_ _2349_ _2350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9020_ _0503_ net29 ci_adder.input_memory\[1\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6428__A1 _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6163_ _1847_ _2240_ _2282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout78_I net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6094_ _2172_ _2214_ _2215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_90_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _1055_ _1225_ _1261_ _1262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4439__B1 _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5045_ _1149_ _1170_ _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7659__B _3459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_36_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6996_ ci_adder.uut_simple_neuron.titan_id_4\[19\] ci_adder.uut_simple_neuron.titan_id_3\[19\]
+ _3086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_67_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8853__CLK net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8804_ _0351_ net17 internal_ih.byte2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5947_ _2068_ _2070_ _2071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_47_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8735_ _0282_ net52 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8666_ ci_adder.stream_o\[18\] ci_adder.output_memory\[18\] _4323_ _4332_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5878_ _1776_ _1878_ _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_75_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7617_ ci_adder.instruction_i\[1\] _3596_ _0704_ _0688_ _3602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_36_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4829_ _0925_ _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__9209__CLK net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8597_ ci_adder.uut_simple_neuron.x0\[27\] ci_adder.input_memory\[1\]\[27\] ci_adder.uut_simple_neuron.x2\[27\]
+ ci_adder.uut_simple_neuron.x3\[27\] _4252_ _4253_ _4289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_105_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7548_ _3540_ _3542_ _3544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7479_ _3486_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4390__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9218_ _0084_ net30 ci_adder.uut_simple_neuron.titan_id_2\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9149_ _0241_ net78 ci_adder.uut_simple_neuron.titan_id_4\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5642__A2 ci_adder.uut_simple_neuron.x3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7919__A1 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8244__I _4052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4381__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8726__CLK net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8876__CLK net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6850_ _2957_ _2958_ _2959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5801_ _1906_ _1927_ _1928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6781_ ci_adder.uut_simple_neuron.x3\[27\] ci_adder.uut_simple_neuron.x3\[28\] _2891_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5732_ _1816_ _1820_ _1860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_91_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8090__S _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8520_ ci_adder.output_memory\[13\] _4212_ _4226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5663_ _1684_ _1792_ _1793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8451_ _4161_ _4170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_115_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5594_ _1711_ _1713_ _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4614_ _0757_ _0777_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7402_ _3422_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8382_ _3654_ _4117_ _4128_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4545_ _0713_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7333_ _3362_ _3363_ _3365_ _3366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_53_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4372__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9003_ _0486_ net65 ci_adder.input_memory\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4476_ _0664_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7264_ ci_adder.uut_simple_neuron.titan_id_1\[4\] ci_adder.uut_simple_neuron.titan_id_0\[4\]
+ _3307_ _3308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_6215_ _2321_ _2333_ _2334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7195_ _3235_ _3236_ _3250_ _3251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6146_ _2178_ _2212_ _2266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6077_ _2098_ ci_adder.uut_simple_neuron.x3\[17\] _2198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6821__A1 _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ _1153_ _1169_ _1177_ _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5927__A3 _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6979_ _3070_ _3071_ _3072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_101_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8718_ _0273_ net71 ci_adder.uut_simple_neuron.x3\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8649_ _3601_ _4323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_106_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5560__A1 _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4363__A2 _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8749__CLK net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5560__B2 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_112_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5863__A2 _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8899__CLK net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_19_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5551__A1 _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5303__A1 ci_adder.uut_simple_neuron.x2\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6000_ _2083_ _2109_ _2121_ _2122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_66_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I spi_cs_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6803__A1 _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7951_ _3866_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ _3007_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7882_ _3824_ _3825_ _3820_ _3821_ _3826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6833_ _2662_ _2664_ _2942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6764_ _2872_ _2873_ _2874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6695_ _2738_ _2741_ _2805_ _2806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5790__A1 ci_adder.uut_simple_neuron.x3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5715_ ci_adder.uut_simple_neuron.x3\[9\] ci_adder.uut_simple_neuron.x3\[10\] _1844_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout7_I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8503_ _0703_ _4212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5646_ _1774_ _1776_ _1777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_8434_ internal_ih.expected_byte_count\[3\] _3958_ _4155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7531__A2 _3524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5577_ _1679_ _1701_ _1710_ _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_5_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8365_ _3616_ _4117_ _4119_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7316_ ci_adder.uut_simple_neuron.titan_id_1\[11\] ci_adder.uut_simple_neuron.titan_id_0\[11\]
+ ci_adder.uut_simple_neuron.titan_id_1\[10\] ci_adder.uut_simple_neuron.titan_id_0\[10\]
+ _3352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8296_ _3645_ _4071_ _4080_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4528_ ci_adder.address_i\[0\] _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_40_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7247_ ci_adder.uut_simple_neuron.titan_id_2\[29\] ci_adder.uut_simple_neuron.titan_id_5\[29\]
+ _3295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4459_ _0655_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7178_ _3235_ _3236_ _3237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6129_ _2098_ _2201_ _2248_ _2249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_99_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A2 ci_adder.uut_simple_neuron.x3\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7770__A2 _3629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9077__CLK net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8914__CLK net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5500_ _1637_ _1639_ _1640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6480_ _2537_ _2540_ _2594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5524__A1 _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5431_ ci_adder.uut_simple_neuron.x2\[25\] ci_adder.uut_simple_neuron.x2\[26\] _1571_
+ _1572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_23_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5362_ _1463_ _1464_ _1504_ _1505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8150_ _3963_ ci_adder.stream_o\[9\] _3981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8313__I1 ci_adder.uut_simple_neuron.x0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7101_ _3169_ _3170_ _3172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8081_ _3934_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7032_ _3113_ _3115_ _3116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5827__A2 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5293_ _1151_ _1436_ _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA_fanout60_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8983_ _0466_ net35 ci_adder.uut_simple_neuron.x0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_77_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7934_ _3680_ ci_adder.uut_simple_neuron.x2\[13\] _3855_ _3858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8529__A1 _4211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7865_ internal_ih.spi_rx_byte_i\[3\] _3805_ _3809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6816_ _1836_ _2851_ _2926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7796_ _3578_ _3749_ _3753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6747_ _2799_ _2857_ _2858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7752__A2 _3629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6678_ _2718_ _2715_ _2789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5629_ _1742_ _1760_ _1761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_61_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8417_ _4146_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_98_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8348_ _3959_ _3965_ _4107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8279_ _4069_ _3838_ _4070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__8607__I2 ci_adder.uut_simple_neuron.x2\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7440__A1 ci_adder.uut_simple_neuron.x0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_1_Left_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_126_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5506__A1 _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5980_ _2094_ _2102_ _2103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4931_ _0807_ _1083_ _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_0_59_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4862_ _1011_ _1016_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7650_ _3611_ _3632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_59_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6601_ _2523_ _2569_ _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_90_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7734__A2 _3659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5745__A1 _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _0948_ _0949_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7581_ _3571_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9320_ _0581_ net47 ci_adder.stream_o\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6532_ _2645_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9242__CLK net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6463_ _2517_ _2577_ _2578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9251_ _0116_ net71 ci_adder.uut_simple_neuron.titan_id_5\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9182_ _0215_ net78 ci_adder.uut_simple_neuron.titan_id_3\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5414_ _1437_ _1539_ _1555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8202_ internal_ih.spi_tx_byte_o\[6\] _3978_ _4028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6394_ _2509_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8133_ _3961_ _3964_ _3965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
XANTENNA__5026__I _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5345_ _0711_ ci_adder.uut_simple_neuron.x2\[27\] _1488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5276_ _1418_ _1420_ _1421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8064_ _3925_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7015_ _3101_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7670__A1 _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8966_ _0449_ net66 ci_adder.uut_simple_neuron.x0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8470__I0 _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7917_ ci_adder.uut_simple_neuron.x2\[5\] _3842_ _3849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8897_ _0044_ net13 ci_adder.value_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7848_ internal_ih.spi_rx_byte_i\[5\] _3787_ _3796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7779_ _3561_ _3562_ _3730_ _3739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_34_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6161__A1 _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7661__A1 ci_adder.value_i\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__A1 internal_ih.byte1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9115__CLK net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4778__A2 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5130_ _1274_ _1277_ _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5061_ _1178_ _1192_ _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8820_ _0367_ net17 internal_ih.byte4\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5966__A1 _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5963_ _1805_ _1917_ _2086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_90_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8751_ _0298_ net65 ci_adder.uut_simple_neuron.x2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4914_ _1064_ _1067_ _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_51_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7702_ _3504_ _3663_ _3675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5894_ _1942_ _1979_ _2019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8682_ _4340_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5718__A1 _1754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4845_ _0969_ _0972_ _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7633_ _1684_ _3617_ _3618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout23_I net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4776_ _0713_ _0900_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8380__A2 _4117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7564_ ci_adder.uut_simple_neuron.x0\[22\] ci_adder.uut_simple_neuron.x0\[23\] _3557_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6515_ _1684_ _1676_ _2455_ _1728_ _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_9303_ _0564_ net45 ci_adder.stream_o\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4941__A2 ci_adder.uut_simple_neuron.x2\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7495_ _3498_ _3499_ _3500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_43_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6446_ _1995_ _2561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_95_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9234_ _0098_ net88 ci_adder.uut_simple_neuron.titan_id_5\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6377_ _1956_ _2433_ _2493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9165_ _0225_ net87 ci_adder.uut_simple_neuron.titan_id_3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8782__CLK net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5328_ _1441_ _1454_ _1471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8116_ _3952_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9096_ _0065_ net48 ci_adder.uut_simple_neuron.titan_id_0\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7643__A1 _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8047_ _3916_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9138__CLK net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5259_ ci_adder.uut_simple_neuron.x2\[24\] ci_adder.uut_simple_neuron.x2\[25\] _1404_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_3_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_82_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5957__A1 _1723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8949_ _0014_ net7 ci_adder.address_i\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9288__CLK net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5709__A1 _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6382__A1 _2491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_91_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4932__A2 ci_adder.uut_simple_neuron.x2\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6134__A1 _2100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4696__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8506__S0 _4206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7634__A1 _3612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4448__A1 internal_ih.byte0\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7810__S _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4999__A2 _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_17_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6373__A1 _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4630_ _0766_ _0769_ _0791_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_72_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6300_ _2414_ _2415_ _2416_ _2417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4561_ _0710_ _0725_ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6125__A1 _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7322__B1 _3354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7280_ _3319_ _3320_ _3321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4492_ internal_ih.byte2\[6\] _0670_ _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6231_ _1907_ _1909_ _2348_ _2349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__8088__S _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6162_ _2279_ _2280_ _2281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6428__A2 _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5113_ _1094_ _1227_ _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__7625__A1 _3608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6093_ _2176_ _2213_ _2214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_90_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5044_ _0870_ _1193_ _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7928__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8803_ _0350_ net17 internal_ih.byte2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6995_ ci_adder.uut_simple_neuron.titan_id_4\[19\] ci_adder.uut_simple_neuron.titan_id_3\[19\]
+ _3085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_48_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5946_ _2017_ _2020_ _2069_ _2070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8734_ spi_interface_cvonk.MOSI_r\[0\] net41 internal_ih.spi_rx_byte_i\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5877_ _1995_ _2001_ _2002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8665_ _4331_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4828_ _0870_ _0983_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7616_ _3600_ _3601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_90_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8596_ ci_adder.output_memory\[27\] _4258_ _4288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4759_ _0892_ _0916_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7547_ _3543_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7478_ _3479_ ci_adder.uut_simple_neuron.x0\[9\] _3485_ _3486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_16_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6429_ _2365_ _2471_ _2544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9217_ _0083_ net30 ci_adder.uut_simple_neuron.titan_id_2\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7864__A1 internal_ih.spi_rx_byte_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9148_ _0240_ net78 ci_adder.uut_simple_neuron.titan_id_4\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9079_ _0532_ net57 ci_adder.output_val_internal\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8416__I0 _3741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4850__A1 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7919__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9303__CLK net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8498__I3 ci_adder.uut_simple_neuron.x3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7855__A1 _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4669__B2 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5800_ _1911_ _1926_ _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6780_ ci_adder.uut_simple_neuron.x3\[26\] _2812_ _2890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8371__S _4122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8583__A2 _4277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5731_ _1790_ _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_85_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5662_ _1681_ _1711_ _1791_ _1792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_45_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8450_ _4165_ _4168_ _4169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5593_ _1725_ _1726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_4613_ _0741_ _0771_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7401_ _3420_ _3421_ _3422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8381_ ci_adder.input_memory\[1\]\[8\] _4118_ _4128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4544_ _0712_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7715__S _3632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7332_ ci_adder.uut_simple_neuron.titan_id_1\[14\] ci_adder.uut_simple_neuron.titan_id_0\[14\]
+ _3365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7846__A1 _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7263_ _3303_ _3305_ _3306_ _3307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6214_ _2332_ _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9002_ _0485_ net66 ci_adder.input_memory\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4475_ internal_ih.byte1\[6\] _0659_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_110_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout90_I net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7194_ ci_adder.uut_simple_neuron.titan_id_2\[19\] ci_adder.uut_simple_neuron.titan_id_5\[19\]
+ _3250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6145_ _2224_ _2264_ _2265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4380__I0 internal_ih.byte4\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6076_ _1999_ _2146_ _2196_ _2197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_99_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8820__CLK net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5027_ _1155_ _1168_ _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5085__A1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6585__A1 _2690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8970__CLK net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6978_ ci_adder.uut_simple_neuron.titan_id_4\[17\] ci_adder.uut_simple_neuron.titan_id_3\[17\]
+ _3071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8717_ _0272_ net71 ci_adder.uut_simple_neuron.x3\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5929_ _1919_ _2052_ _2053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_101_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6337__A1 _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8648_ _4322_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8579_ ci_adder.output_val_internal\[23\] _4249_ _4275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4899__A1 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7837__A1 _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8637__I0 ci_adder.stream_o\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5551__A2 ci_adder.uut_simple_neuron.x3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5303__A2 ci_adder.uut_simple_neuron.x2\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7950_ _3723_ _1233_ _3855_ _3866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8993__CLK net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6901_ ci_adder.uut_simple_neuron.titan_id_4\[4\] ci_adder.uut_simple_neuron.titan_id_3\[4\]
+ _3006_ _3007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_7881_ _3818_ _3825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6832_ _2662_ _2664_ _2941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6763_ _2797_ _2858_ _2873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_18_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6694_ _2742_ _2746_ _2805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5714_ ci_adder.uut_simple_neuron.x3\[7\] _1804_ _1842_ _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_85_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8502_ _4161_ _4211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5645_ ci_adder.uut_simple_neuron.x3\[6\] _1775_ _1776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_8433_ _0583_ _3958_ _4154_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5576_ ci_adder.uut_simple_neuron.x3\[3\] ci_adder.uut_simple_neuron.x3\[4\] _1710_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8364_ ci_adder.input_memory\[1\]\[0\] _4118_ _4119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7315_ _3342_ _3347_ _3351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8295_ _3469_ _4072_ _4080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4527_ ci_adder.address_i\[1\] _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7246_ ci_adder.uut_simple_neuron.titan_id_2\[29\] ci_adder.uut_simple_neuron.titan_id_5\[29\]
+ _3294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4458_ internal_ih.byte0\[6\] _0648_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7177_ ci_adder.uut_simple_neuron.titan_id_2\[19\] ci_adder.uut_simple_neuron.titan_id_5\[19\]
+ _3236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6128_ ci_adder.uut_simple_neuron.x3\[17\] _2200_ _2248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4389_ internal_ih.byte4\[7\] internal_ih.byte3\[7\] _0599_ _0617_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4817__B ci_adder.uut_simple_neuron.x2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6059_ _1772_ _2136_ _2180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8547__A2 _4247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8716__CLK net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8866__CLK net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6797__A1 _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8538__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6549__A1 _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7210__A2 ci_adder.uut_simple_neuron.titan_id_5\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5430_ _1348_ _1445_ _1571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6721__A1 _1807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5361_ _1460_ _1462_ _1504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5292_ _1084_ _1435_ _1436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8080_ internal_ih.byte6\[3\] internal_ih.byte5\[3\] _3930_ _3934_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8474__A1 ci_adder.output_memory\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7100_ _3171_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7031_ _3110_ _3111_ _3114_ _3115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8096__S _3825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8982_ _0465_ net26 ci_adder.uut_simple_neuron.x0\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_117_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9171__CLK net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7933_ _3857_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout53_I net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5460__A1 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7864_ internal_ih.spi_rx_byte_i\[1\] internal_ih.spi_rx_byte_i\[0\] internal_ih.spi_rx_byte_i\[2\]
+ _3808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_6815_ _1841_ _1851_ _2925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7795_ _2953_ _3612_ _3752_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7201__A2 ci_adder.uut_simple_neuron.titan_id_5\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6746_ _2842_ _2856_ _2857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_61_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6677_ _2706_ _2786_ _2788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5628_ _1745_ _1759_ _1760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7760__I0 _3723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8416_ _3741_ ci_adder.input_memory\[1\]\[25\] _4139_ _4146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5559_ _1684_ _1676_ _1679_ _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_13_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8347_ _4106_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8278_ _3608_ _3609_ _4069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7229_ _3277_ _3279_ _3280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8607__I3 ci_adder.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7440__A2 _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A1 _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9044__CLK net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8456__A1 _4165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_102_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8208__A1 _3811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4930_ _1079_ _1082_ _0963_ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_4
XANTENNA__8443__I _4161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_111_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4861_ _1012_ _1015_ _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
X_6600_ _2712_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5745__A2 _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4792_ _0919_ _0920_ _0947_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_55_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7580_ _3569_ _3570_ _3571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6531_ _2581_ _2644_ _2645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_55_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6462_ _2576_ _2577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7742__I0 _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9250_ _0115_ net71 ci_adder.uut_simple_neuron.titan_id_5\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6393_ _2504_ _2505_ _2508_ _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_9181_ _0214_ net77 ci_adder.uut_simple_neuron.titan_id_3\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5413_ _1521_ _1538_ _1554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8201_ ci_adder.stream_o\[30\] _3959_ _4026_ _4027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_120_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5344_ _1484_ _1486_ _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7723__S _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8132_ internal_ih.data_pointer\[0\] _3964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5275_ _1419_ _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8063_ internal_ih.byte5\[3\] internal_ih.byte4\[3\] _3919_ _3925_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7014_ _3099_ _3100_ _3101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5433__A1 ci_adder.uut_simple_neuron.x2\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8965_ _0448_ net66 ci_adder.uut_simple_neuron.x0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7916_ _3636_ _3841_ _3848_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_54_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8896_ _0033_ net13 ci_adder.value_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7847_ internal_ih.spi_tx_byte_o\[4\] _3779_ _3784_ internal_ih.spi_rx_byte_i\[4\]
+ _3795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7981__I0 internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7778_ ci_adder.value_i\[25\] _3659_ _3738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6729_ _2833_ _2839_ _2840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__9067__CLK net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8904__CLK net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7661__A2 _3619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6048__I _2169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5672__A1 ci_adder.uut_simple_neuron.x3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__A2 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4778__A3 ci_adder.uut_simple_neuron.x2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8516__I2 _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5060_ _1209_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5663__A1 _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8601__A1 ci_adder.output_memory\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5962_ _2042_ _2059_ _2084_ _2085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_84_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8750_ _0297_ net52 internal_ih.received_byte_count\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4913_ _0996_ _1065_ _1066_ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7701_ ci_adder.value_i\[12\] _3659_ _3674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5893_ _1942_ _1979_ _2018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_90_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8681_ ci_adder.stream_o\[25\] ci_adder.output_memory\[25\] _4334_ _4340_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4844_ _0955_ _0997_ _0998_ _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7632_ _3611_ _3617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__8460__S0 _4166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4775_ _0894_ _0931_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4777__I0 ci_adder.uut_simple_neuron.x2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout16_I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7563_ ci_adder.uut_simple_neuron.x0\[23\] ci_adder.uut_simple_neuron.x0\[24\] _3556_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6514_ _2588_ _2627_ _2628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9302_ _0563_ net45 ci_adder.stream_o\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9233_ _0097_ net85 ci_adder.uut_simple_neuron.titan_id_5\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7494_ _3487_ _3493_ _3494_ _3499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_15_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6445_ _2558_ _2559_ _2560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_95_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8927__CLK net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6376_ _1962_ _2432_ _2492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9164_ _0224_ net85 ci_adder.uut_simple_neuron.titan_id_3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5327_ _1468_ _1469_ _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_11_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8115_ internal_ih.current_instruction\[4\] _3947_ _3952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_9095_ ci_adder.uut_simple_neuron.x0\[0\] net48 ci_adder.uut_simple_neuron.titan_id_0\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7643__A2 _3617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8046_ internal_ih.byte4\[3\] internal_ih.byte3\[3\] _3908_ _3916_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5258_ ci_adder.uut_simple_neuron.x2\[24\] ci_adder.uut_simple_neuron.x2\[25\] _1403_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_3_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5189_ _1110_ _1333_ _1334_ _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8948_ _0013_ net7 ci_adder.address_i\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5957__A2 _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8879_ _0426_ net56 ci_adder.output_memory\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5709__A2 _1807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7954__I0 _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7882__A2 _3825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8506__S1 _4207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5645__A1 ci_adder.uut_simple_neuron.x3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7634__A2 _3616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6070__A1 _1807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4560_ _0722_ _0723_ _0726_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4384__B2 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4491_ _0672_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6230_ _1948_ _1923_ _2348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5884__A1 _1947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6161_ _0162_ _2232_ _2280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5112_ _1091_ _1259_ _1016_ _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6092_ _2178_ _2212_ _2213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5636__A1 _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4439__A2 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5043_ _1178_ _1192_ _1193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_33_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8802_ _0349_ net23 internal_ih.byte2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6994_ _3084_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_36_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5945_ _1981_ _2016_ _2069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_88_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8733_ net3 net41 spi_interface_cvonk.MOSI_r\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5876_ _1880_ _2000_ _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8664_ ci_adder.stream_o\[17\] ci_adder.output_memory\[17\] _4323_ _4331_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4827_ _0953_ _0982_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7615_ ci_adder.instruction_i\[0\] ci_adder.instruction_i\[1\] ci_adder.stream_enabled
+ _3596_ _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_29_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7561__A1 ci_adder.uut_simple_neuron.x0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8595_ _4257_ _4284_ _4286_ _4287_ _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4758_ _0804_ _0915_ _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7546_ _3540_ _3542_ _3543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4375__B2 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4689_ _0811_ _0834_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7477_ _3484_ _3481_ _3485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6428_ _2365_ _2471_ _2543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9216_ _0082_ net30 ci_adder.uut_simple_neuron.titan_id_2\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7864__A2 internal_ih.spi_rx_byte_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9147_ _0239_ net78 ci_adder.uut_simple_neuron.titan_id_4\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5875__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6359_ _2471_ _2474_ _2475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8113__I0 internal_ih.spi_rx_byte_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5627__A1 _1723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8664__I1 ci_adder.output_memory\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9078_ _0531_ net55 ci_adder.output_val_internal\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9255__CLK net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8029_ internal_ih.byte3\[3\] internal_ih.byte2\[3\] _3897_ _3907_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5866__A1 _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6291__A1 _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8652__S _4323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ _1858_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8451__I _4161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5661_ _1686_ _1769_ _1791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7400_ ci_adder.uut_simple_neuron.titan_id_1\[27\] ci_adder.uut_simple_neuron.titan_id_0\[27\]
+ _3421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5592_ _1723_ _1724_ _1725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__9128__CLK net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4612_ _0765_ _0775_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8380_ _3650_ _4117_ _4127_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ _0711_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7331_ _3364_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7262_ ci_adder.uut_simple_neuron.titan_id_1\[3\] ci_adder.uut_simple_neuron.titan_id_0\[3\]
+ _3306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6213_ _2328_ _2331_ _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5857__A1 _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9001_ _0484_ net66 ci_adder.input_memory\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4474_ _0663_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7193_ _3241_ _3246_ _3249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6144_ _2226_ _2263_ _2264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6075_ _2143_ _2195_ _2196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5026_ _1176_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_49_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6977_ _3068_ _3069_ _3070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5928_ _2049_ _2051_ _2052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8716_ _0271_ net72 ci_adder.uut_simple_neuron.x3\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_101_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5859_ _1982_ _1983_ _1984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8647_ ci_adder.stream_o\[9\] ci_adder.output_memory\[9\] _4312_ _4322_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8578_ _4260_ _4273_ _4274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7529_ _3528_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8334__I0 _3741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4371__I1 internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8637__I1 ci_adder.output_memory\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6025__A1 _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6005__B _2126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7525__A1 ci_adder.uut_simple_neuron.x0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5839__A1 _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5303__A3 ci_adder.uut_simple_neuron.x2\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8446__I _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6900_ _3002_ _3004_ _3005_ _3006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7880_ _3807_ _3808_ _3814_ _3824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6831_ _2872_ _2873_ _2936_ _2940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_46_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4578__A1 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6762_ _2799_ _2871_ _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8501_ _4162_ _4205_ _4209_ _4210_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6693_ _2802_ _2752_ _2803_ _2804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5713_ ci_adder.uut_simple_neuron.x3\[8\] ci_adder.uut_simple_neuron.x3\[9\] _1842_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7516__A1 ci_adder.uut_simple_neuron.x0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5644_ ci_adder.uut_simple_neuron.x3\[7\] ci_adder.uut_simple_neuron.x3\[8\] _1775_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_73_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8432_ internal_ih.spi_rx_byte_i\[1\] internal_ih.spi_rx_byte_i\[2\] _3958_ _4154_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_33_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8363_ _4116_ _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5575_ _1677_ _1703_ _1708_ _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7314_ _3329_ _3338_ _3349_ _3350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_13_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8294_ _3641_ _4071_ _4079_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4526_ ci_adder.address_i\[22\] ci_adder.address_i\[23\] _0690_ _0695_ _0696_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_13_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4457_ _0654_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7245_ _3293_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7176_ _3231_ _3232_ _3234_ _3235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6127_ _2051_ _2203_ _2246_ _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4388_ _0616_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6058_ _1778_ _2135_ _2179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5009_ ci_adder.uut_simple_neuron.x2\[18\] ci_adder.uut_simple_neuron.x2\[19\] _1160_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4569__A1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7755__A1 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8307__I0 _3677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_15_Left_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_115_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6494__A1 _2249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6246__A1 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_24_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_125_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8810__CLK net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_33_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5360_ _1500_ _1502_ _1503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_77_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5291_ _1302_ _1303_ _1399_ _1434_ _1311_ _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_11_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7030_ ci_adder.uut_simple_neuron.titan_id_4\[25\] ci_adder.uut_simple_neuron.titan_id_3\[25\]
+ _3114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6485__A1 _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6237__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9316__CLK net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8981_ _0464_ net33 ci_adder.uut_simple_neuron.x0\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4799__A1 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7932_ _3677_ _0899_ _3855_ _3857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7863_ _3804_ internal_ih.spi_rx_byte_i\[3\] _3806_ _3807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_4
XANTENNA_fanout46_I net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6814_ _2922_ _2923_ _2924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7794_ _3632_ _3751_ _3752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6745_ _2844_ _2855_ _2856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4971__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6676_ _2787_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8415_ _4145_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5627_ _1723_ _1748_ _1758_ _1759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_103_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7760__I1 _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5558_ _1675_ _1693_ _1694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8346_ _3768_ ci_adder.uut_simple_neuron.x0\[31\] _4070_ _4106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8277_ _0587_ _3820_ _3822_ _3958_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4509_ _0681_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5489_ _1560_ _1605_ _1628_ _1629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7228_ _3274_ _3275_ _3278_ _3279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6228__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7159_ ci_adder.uut_simple_neuron.titan_id_2\[16\] ci_adder.uut_simple_neuron.titan_id_5\[16\]
+ _3221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_29_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7728__A1 _3619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6400__A1 _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8833__CLK net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4962__A1 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7900__A1 _3826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4714__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4860_ _1013_ _1014_ _0894_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_28_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8660__S _4323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6530_ _2582_ _2643_ _2644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4791_ _0919_ _0920_ _0947_ _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7990__I1 internal_ih.byte0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6461_ _2518_ _2575_ _2576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6392_ _2506_ _2507_ _2508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9180_ _0213_ net79 ci_adder.uut_simple_neuron.titan_id_3\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5412_ _1551_ _1552_ _1553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7742__I1 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8200_ _3960_ _4023_ _4025_ _3815_ _4026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5343_ _1485_ _1403_ _1486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8131_ _3962_ _3963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_112_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5274_ _1385_ _1386_ _1417_ _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_11_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8062_ _3924_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7013_ ci_adder.uut_simple_neuron.titan_id_4\[23\] ci_adder.uut_simple_neuron.titan_id_3\[23\]
+ _3100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8470__I2 ci_adder.uut_simple_neuron.x2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8964_ _0447_ net56 ci_adder.uut_simple_neuron.x0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_7915_ ci_adder.uut_simple_neuron.x2\[4\] _3842_ _3848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8895_ _0442_ net18 ci_adder.output_memory\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_54_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7846_ _3770_ _3793_ _3794_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7186__A2 ci_adder.uut_simple_neuron.titan_id_5\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4989_ _1139_ _1140_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7777_ _3737_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6728_ _2836_ _2838_ _2839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6659_ _1770_ _1772_ _2771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8329_ _3728_ _4072_ _4097_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5121__A1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5672__A2 ci_adder.uut_simple_neuron.x3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6621__A1 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4778__A4 _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5188__A1 _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8374__A1 _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9011__CLK net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8516__I3 ci_adder.uut_simple_neuron.x3\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9161__CLK net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8729__CLK net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5143__I _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8879__CLK net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ _2045_ _2058_ _2084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4912_ _0999_ _1024_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7700_ _3673_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8680_ _4339_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5892_ _1981_ _2016_ _2017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_90_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8365__A1 _3616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7631_ ci_adder.value_i\[0\] _3613_ _3615_ _3616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_118_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4843_ _0959_ _0981_ _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8460__S1 _4167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4774_ _0899_ ci_adder.uut_simple_neuron.x2\[13\] _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4926__A1 _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7562_ _3555_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6513_ _2616_ _2626_ _2627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7493_ _3487_ _3493_ _3489_ _3490_ _3488_ _3498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_9301_ _0562_ net46 ci_adder.stream_o\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6444_ _1715_ _2495_ _2559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9232_ _0126_ net85 ci_adder.uut_simple_neuron.titan_id_5\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7715__I1 ci_adder.uut_simple_neuron.x3\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6375_ _2489_ _2490_ _2491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9163_ _0223_ net85 ci_adder.uut_simple_neuron.titan_id_3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5326_ _1151_ _1436_ _1469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8114_ _3951_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9094_ _0547_ net45 ci_adder.output_val_internal\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5103__A1 _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5257_ _1353_ _1399_ _1402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8045_ _3915_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5188_ _1151_ _1319_ _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7651__I0 _3631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8947_ _0011_ net7 ci_adder.address_i\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8878_ _0425_ net48 ci_adder.output_memory\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7954__I1 ci_adder.uut_simple_neuron.x2\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7829_ spi_interface_cvonk.state\[1\] spi_interface_cvonk.state\[0\] _3781_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_93_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5590__A1 _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_7_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4384__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4490_ internal_ih.byte2\[5\] _0670_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_122_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6160_ _1836_ _1851_ _2279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5111_ _1094_ _1227_ _1259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_0_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6091_ _2185_ _2211_ _2212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5636__A2 _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5042_ _1156_ _1191_ _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9057__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8801_ _0348_ net23 internal_ih.byte2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8586__A1 ci_adder.output_memory\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6993_ ci_adder.uut_simple_neuron.titan_id_4\[19\] ci_adder.uut_simple_neuron.titan_id_3\[19\]
+ _3083_ _3084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_88_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7729__S _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5944_ _2066_ _2067_ _2068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8732_ spi_interface_cvonk.SS_r\[1\] net52 spi_interface_cvonk.SS_r\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5875_ _1997_ _1999_ _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_48_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8663_ _4330_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4826_ _0955_ _0959_ _0981_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__7936__I1 ci_adder.uut_simple_neuron.x2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7614_ _3598_ _3599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8594_ ci_adder.output_val_internal\[26\] _4249_ _4287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7545_ _3524_ ci_adder.uut_simple_neuron.x0\[18\] _3532_ _3534_ _3541_ _3542_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_16_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4375__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4757_ _0879_ _0914_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4688_ _0836_ _0837_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7476_ _3470_ _3479_ _3484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8510__A1 ci_adder.output_memory\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6427_ _2418_ _2541_ _2542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9215_ _0081_ net30 ci_adder.uut_simple_neuron.titan_id_2\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9146_ _0238_ net78 ci_adder.uut_simple_neuron.titan_id_4\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5875__A2 _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6358_ ci_adder.uut_simple_neuron.x3\[23\] _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_3_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ _1444_ _1452_ _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6289_ _2404_ _2356_ _2405_ _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9077_ _0530_ net54 ci_adder.output_val_internal\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8028_ _3906_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8329__A1 _3728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7552__A2 ci_adder.uut_simple_neuron.x0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5563__A1 _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6815__A1 _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8917__CLK net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ _1785_ _1787_ _1790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_45_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4611_ _0770_ _0771_ _0774_ _0742_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5591_ _1675_ _1689_ _1724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4542_ ci_adder.uut_simple_neuron.x2\[1\] _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7330_ _3362_ _3363_ _3364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_52_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5306__A1 _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4473_ internal_ih.byte1\[5\] _0659_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7261_ ci_adder.uut_simple_neuron.titan_id_1\[3\] ci_adder.uut_simple_neuron.titan_id_0\[3\]
+ _3305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6212_ _2066_ _2072_ _2330_ _2331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5857__A2 _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9000_ _0483_ net58 ci_adder.input_memory\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7192_ ci_adder.uut_simple_neuron.titan_id_2\[21\] ci_adder.uut_simple_neuron.titan_id_5\[21\]
+ _3248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6143_ _2235_ _2262_ _2263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_fanout76_I net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6074_ _2050_ _2144_ _2195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5025_ _1173_ _1175_ _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_49_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6976_ _3065_ _3066_ _3069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5793__A1 _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5927_ ci_adder.uut_simple_neuron.x3\[13\] ci_adder.uut_simple_neuron.x3\[14\] _2050_
+ _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_8715_ _0270_ net73 ci_adder.uut_simple_neuron.x3\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_101_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5858_ _1721_ _1951_ _1983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8646_ _4321_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5545__A1 _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5789_ ci_adder.uut_simple_neuron.x3\[10\] ci_adder.uut_simple_neuron.x3\[11\] _1916_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4809_ _0963_ _0940_ _0964_ _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8577_ ci_adder.uut_simple_neuron.x0\[23\] ci_adder.input_memory\[1\]\[23\] ci_adder.uut_simple_neuron.x2\[23\]
+ _2474_ _4252_ _4253_ _4273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_44_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7528_ ci_adder.uut_simple_neuron.x0\[16\] _3524_ _3527_ _3528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7459_ ci_adder.uut_simple_neuron.x0\[6\] _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__9222__CLK net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_79_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9129_ _0163_ net88 ci_adder.uut_simple_neuron.titan_id_4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_19_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_88_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8552__I _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5784__A1 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_97_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7787__B _3745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6830_ _2939_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6761_ _2857_ _2871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5712_ _1732_ _1806_ _1840_ _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_85_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8013__I0 internal_ih.byte2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8500_ ci_adder.output_val_internal\[9\] _4203_ _4210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6692_ _2731_ _2747_ _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9245__CLK net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5643_ ci_adder.uut_simple_neuron.x3\[5\] _1753_ _1773_ _1774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_73_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8431_ _4153_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5574_ _1700_ _1702_ _1708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_14_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8362_ _4116_ _4117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_115_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7313_ _3337_ _3340_ _3349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4525_ _0691_ _0692_ _0693_ _0694_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_13_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7742__S _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8572__S0 _4252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8293_ _3459_ _4072_ _4079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7244_ ci_adder.uut_simple_neuron.titan_id_2\[29\] ci_adder.uut_simple_neuron.titan_id_5\[29\]
+ _3292_ _3293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_1_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4456_ internal_ih.byte0\[5\] _0648_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7175_ ci_adder.uut_simple_neuron.titan_id_2\[18\] ci_adder.uut_simple_neuron.titan_id_5\[18\]
+ _3234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4387_ internal_ih.byte7\[6\] _0603_ _0615_ net14 _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6126_ _2199_ _2245_ _2246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6057_ _2130_ _2154_ _2177_ _2178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5008_ _1012_ _1015_ _1090_ _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_68_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7755__A2 _3612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6959_ ci_adder.uut_simple_neuron.titan_id_4\[13\] ci_adder.uut_simple_neuron.titan_id_3\[13\]
+ _3055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4569__A2 _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8004__I0 internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8629_ ci_adder.stream_o\[0\] ci_adder.output_memory\[0\] _4312_ _4313_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7691__A1 _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_73_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7746__A2 _3659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9268__CLK net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6182__A1 _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8658__S _4323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5290_ _1310_ _1399_ _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8554__S0 _4252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7682__A1 _3479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4496__A1 internal_ih.byte3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8393__S _4122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8980_ _0463_ net33 ci_adder.uut_simple_neuron.x0\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_78_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7931_ _3856_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7862_ internal_ih.spi_rx_byte_i\[1\] internal_ih.spi_rx_byte_i\[0\] _3805_ _3806_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6813_ _2833_ _2839_ _2923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5748__A1 _1754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout39_I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7793_ _3748_ _3750_ _3751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6744_ _2847_ _2854_ _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_92_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ _2717_ _2786_ _2787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5626_ _1750_ _1756_ _1757_ _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_60_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8414_ _3736_ ci_adder.input_memory\[1\]\[24\] _4139_ _4145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6173__A1 _1958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5557_ _1690_ _1692_ _1693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_5_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8345_ _4105_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5488_ _1525_ _1627_ _1628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4508_ internal_ih.byte3\[6\] _0597_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8276_ _4068_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7673__A1 ci_adder.uut_simple_neuron.x3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7227_ ci_adder.uut_simple_neuron.titan_id_2\[26\] ci_adder.uut_simple_neuron.titan_id_5\[26\]
+ _3278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4439_ internal_ih.byte6\[5\] _0635_ _0619_ internal_ih.byte2\[5\] _0645_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7158_ _3216_ _3218_ _3219_ _3220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6109_ _1807_ _2190_ _2229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7089_ _3160_ _3161_ _3162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_29_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5739__A1 _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6400__A2 _2072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6164__A1 _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8536__S0 _4206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7664__A1 _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4650__A1 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4790_ _0922_ _0946_ _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_86_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6460_ _2571_ _2574_ _2575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6391_ _2381_ _2379_ _2441_ _2507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5902__A1 _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5411_ _1470_ _1541_ _1552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5342_ ci_adder.uut_simple_neuron.x2\[26\] _1485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8130_ _3961_ _3962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_11_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8061_ internal_ih.byte5\[2\] internal_ih.byte4\[2\] _3919_ _3924_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7655__A1 _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7012_ _3095_ _3097_ _3098_ _3099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_5273_ _1385_ _1386_ _1417_ _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4469__A1 internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8470__I3 ci_adder.uut_simple_neuron.x3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8963_ _0446_ net61 ci_adder.uut_simple_neuron.x0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_7914_ _3847_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8894_ _0441_ net22 ci_adder.output_memory\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_54_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7845_ internal_ih.spi_rx_byte_i\[4\] _3787_ _3794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4988_ _1072_ _1102_ _1104_ _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7776_ _3736_ _2538_ _3692_ _3737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6727_ _1847_ _2837_ _2838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6658_ _2768_ _2769_ _2770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5609_ _1741_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6589_ _2586_ _2639_ _2702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8328_ ci_adder.uut_simple_neuron.x0\[22\] _4076_ _4097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7646__A1 ci_adder.uut_simple_neuron.x0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7930__S _3855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8259_ ci_adder.uut_simple_neuron.titan_id_6\[23\] _4060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_6_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8800__CLK net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8374__A2 _4117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8950__CLK net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6137__A1 _1958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9306__CLK net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6688__A2 _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7904__I _3840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_70_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4871__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5960_ _2079_ _2082_ _2083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5891_ _2011_ _2015_ _2016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4911_ _0999_ _1024_ _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_51_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8365__A2 _4117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7630_ ci_adder.uut_simple_neuron.x0\[0\] _3614_ _3615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6376__A1 _1962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4842_ _0959_ _0981_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4773_ _0715_ _0928_ _0902_ _0929_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7561_ ci_adder.uut_simple_neuron.x0\[22\] ci_adder.uut_simple_neuron.x0\[23\] _3554_
+ _3555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_7_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8117__A2 _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6512_ _2619_ _2625_ _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6128__A1 ci_adder.uut_simple_neuron.x3\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7492_ ci_adder.uut_simple_neuron.x0\[11\] ci_adder.uut_simple_neuron.x0\[12\] _3497_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_15_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9300_ _0561_ net46 ci_adder.stream_o\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6443_ _1989_ _2004_ _2558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9231_ _0125_ net86 ci_adder.uut_simple_neuron.titan_id_5\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7876__A1 _3811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6374_ _1704_ _2407_ _2490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9162_ _0200_ net85 ci_adder.uut_simple_neuron.titan_id_3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5325_ _1084_ _1435_ _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8113_ internal_ih.spi_rx_byte_i\[3\] internal_ih.current_instruction\[3\] _3947_
+ _3951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9093_ _0546_ net54 ci_adder.output_val_internal\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5256_ _1351_ _1353_ _1354_ _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__8823__CLK net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8044_ internal_ih.byte4\[2\] internal_ih.byte3\[2\] _3908_ _3915_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6851__A2 _2956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5187_ _1304_ _1333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4862__A1 _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7651__I1 ci_adder.uut_simple_neuron.x3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8973__CLK net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8946_ _0010_ net7 ci_adder.address_i\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8877_ _0424_ net63 ci_adder.output_memory\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_104_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7828_ spi_interface_cvonk.SCLK_r\[2\] _3771_ _3780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__9128__D _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8108__A2 _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7759_ _3619_ _3720_ _3721_ _3722_ _3723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_117_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6119__A1 _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7925__S _3846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8292__A1 _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7095__A2 ci_adder.uut_simple_neuron.titan_id_5\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4853__A1 _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4369__B1 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8846__CLK net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8666__S _4323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6090_ _2188_ _2210_ _2211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_85_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5110_ _1232_ _1236_ _1257_ _1233_ _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__8283__A1 _3616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5041_ _1180_ _1190_ _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8996__CLK net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_108_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8800_ _0347_ net19 internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6992_ _3073_ _3078_ _3079_ _3081_ _3082_ _3083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_8731_ spi_interface_cvonk.SS_r\[0\] net52 spi_interface_cvonk.SS_r\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5943_ _2011_ _2022_ _2065_ _2067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5874_ ci_adder.uut_simple_neuron.x3\[12\] _1998_ _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_47_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8662_ ci_adder.stream_o\[16\] ci_adder.output_memory\[16\] _4323_ _4330_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5021__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4825_ _0969_ _0972_ _0980_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_63_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout21_I net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7613_ _0700_ _3597_ _3598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8593_ _4260_ _4285_ _4286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_117_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7544_ _3535_ _3541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_50_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4756_ _0893_ _0913_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7849__A1 _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4687_ _0832_ _0839_ _0846_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7475_ _3483_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8510__A2 _4212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6521__A1 _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6426_ _2537_ _2540_ _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9214_ _0080_ net38 ci_adder.uut_simple_neuron.titan_id_2\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9145_ _0237_ net79 ci_adder.uut_simple_neuron.titan_id_4\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6357_ ci_adder.uut_simple_neuron.x3\[20\] _2423_ _2472_ _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4383__I0 internal_ih.byte4\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5308_ _1402_ _1451_ _1452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_126_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6288_ _1921_ _2355_ _2405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9001__CLK net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9076_ _0529_ net54 ci_adder.output_val_internal\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5239_ _1384_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8027_ internal_ih.byte3\[2\] internal_ih.byte2\[2\] _3897_ _3906_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7624__I1 _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9151__CLK net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5260__A1 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8329__A2 _4072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8929_ _0012_ net8 ci_adder.address_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8869__CLK net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8568__A2 _4265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5251__A1 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7629__I _3599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8040__I1 internal_ih.byte3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4610_ _0773_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6751__A1 _2720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5590_ _1684_ _1690_ _1723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_25_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7792__C _3599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4541_ _0709_ _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_53_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4472_ _0662_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7260_ _3304_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6211_ _2323_ _2329_ _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9024__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7191_ _3247_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6142_ _2238_ _2261_ _2262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6073_ _2148_ _2151_ _2193_ _2194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4817__A1 _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5024_ _1138_ _1143_ _1174_ _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9174__CLK net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout69_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6975_ ci_adder.uut_simple_neuron.titan_id_4\[16\] ci_adder.uut_simple_neuron.titan_id_3\[16\]
+ _3068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5793__A2 _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5926_ ci_adder.uut_simple_neuron.x3\[15\] _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8714_ _0269_ net73 ci_adder.uut_simple_neuron.x3\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8645_ ci_adder.stream_o\[8\] ci_adder.output_memory\[8\] _4312_ _4321_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5857_ _1704_ _1950_ _1982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8582__I2 ci_adder.uut_simple_neuron.x2\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5788_ _1776_ _1881_ _1914_ _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_91_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4808_ _0928_ _0909_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8576_ ci_adder.output_memory\[23\] _4258_ _4272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4739_ _0834_ _0852_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7527_ _3525_ _3526_ _3527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7458_ _3468_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8495__A1 ci_adder.output_memory\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6409_ _2494_ _2496_ _2524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7389_ ci_adder.uut_simple_neuron.titan_id_1\[25\] ci_adder.uut_simple_neuron.titan_id_0\[25\]
+ _3412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_40_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9128_ _0162_ net88 ci_adder.uut_simple_neuron.titan_id_4\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9059_ ci_adder.input_memory\[1\]\[27\] net31 ci_adder.uut_simple_neuron.titan_id_1\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_67_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6981__A1 ci_adder.uut_simple_neuron.titan_id_4\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6733__A1 _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9047__CLK net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8486__A1 _4165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7912__I _3840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9197__CLK net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8410__A1 ci_adder.input_memory\[1\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6760_ _2859_ _2863_ _2870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5711_ _1803_ _1805_ _1840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6972__A1 ci_adder.uut_simple_neuron.titan_id_4\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8013__I1 internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6691_ _2731_ _2747_ _2802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5642_ ci_adder.uut_simple_neuron.x3\[6\] ci_adder.uut_simple_neuron.x3\[7\] _1773_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7772__I0 _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8430_ _3976_ internal_ih.expected_byte_count\[0\] _3958_ _4153_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5573_ _1707_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8361_ _3607_ _4069_ _4116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_41_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7312_ _3348_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4524_ ci_adder.address_i\[9\] ci_adder.address_i\[8\] ci_adder.address_i\[7\] ci_adder.address_i\[6\]
+ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_13_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8477__A1 ci_adder.output_val_internal\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8292_ _3636_ _4071_ _4078_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7243_ _3288_ _3290_ _3291_ _3292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8572__S1 _4253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4455_ _0653_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7174_ _3233_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4386_ internal_ih.byte4\[6\] internal_ih.byte3\[6\] _0599_ _0615_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6125_ _2098_ _2201_ _2245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5342__I ci_adder.uut_simple_neuron.x2\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6056_ _2133_ _2153_ _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5007_ _1095_ _1125_ _1127_ _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_68_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7204__A2 ci_adder.uut_simple_neuron.titan_id_5\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6958_ _3054_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5909_ _2032_ _2033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6889_ _2997_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8004__I1 internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8628_ _3601_ _4312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_24_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8559_ _0703_ _4258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_122_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8907__CLK net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5454__A1 _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5206__A1 ci_adder.uut_simple_neuron.x2\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8546__I2 ci_adder.uut_simple_neuron.x2\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6182__A2 ci_adder.uut_simple_neuron.x3\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8459__A1 ci_adder.output_memory\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8554__S1 _4253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7798__B _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7930_ _3672_ ci_adder.uut_simple_neuron.x2\[11\] _3855_ _3856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7861_ internal_ih.spi_rx_byte_i\[7\] internal_ih.spi_rx_byte_i\[6\] internal_ih.spi_rx_byte_i\[5\]
+ internal_ih.spi_rx_byte_i\[4\] _3805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6812_ _2836_ _2838_ _2922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9212__CLK net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8490__S0 _4166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7792_ _3578_ _3749_ _3744_ ci_adder.uut_simple_neuron.x0\[27\] _3599_ _3750_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_6743_ _0162_ _2853_ _2854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6674_ _2718_ _2785_ _2786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_18_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5625_ _0162_ _1700_ _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_8413_ _4144_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_21_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5556_ ci_adder.uut_simple_neuron.x3\[1\] _1691_ _1692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_4
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8344_ _3765_ ci_adder.uut_simple_neuron.x0\[30\] _4070_ _4105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5487_ _1608_ _1626_ _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4507_ _0680_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8275_ ci_adder.uut_simple_neuron.titan_id_6\[31\] _4068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7673__A2 _3617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7226_ ci_adder.uut_simple_neuron.titan_id_2\[27\] ci_adder.uut_simple_neuron.titan_id_5\[27\]
+ _3277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4438_ _0644_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7157_ ci_adder.uut_simple_neuron.titan_id_2\[15\] ci_adder.uut_simple_neuron.titan_id_5\[15\]
+ _3219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4369_ net14 _0600_ _0603_ internal_ih.byte7\[0\] _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6108_ _1684_ _2182_ _2227_ _2228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7088_ _3157_ _3158_ _3161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6039_ _2112_ _2114_ _2161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_69_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5739__A2 _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4411__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7736__I0 _3703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8536__S1 _4207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8558__I _4161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5675__A1 ci_adder.uut_simple_neuron.x3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8613__A1 _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5978__A2 _2100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4650__A2 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7975__I0 internal_ih.byte0\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6390_ _2442_ _2447_ _2506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5410_ _1518_ _1540_ _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5341_ ci_adder.uut_simple_neuron.x2\[24\] ci_adder.uut_simple_neuron.x2\[25\] ci_adder.uut_simple_neuron.x2\[26\]
+ _1484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8060_ _3923_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7011_ ci_adder.uut_simple_neuron.titan_id_4\[22\] ci_adder.uut_simple_neuron.titan_id_3\[22\]
+ _3098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5272_ _0994_ _1416_ _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4469__A2 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5418__A1 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8962_ _0445_ net56 ci_adder.uut_simple_neuron.x0\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_7913_ _3631_ _0722_ _3846_ _3847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout51_I net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7748__S _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8893_ _0440_ net32 ci_adder.output_memory\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7844_ internal_ih.spi_tx_byte_o\[3\] _3779_ _3784_ internal_ih.spi_rx_byte_i\[3\]
+ _3793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_65_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7775_ ci_adder.value_i\[24\] _3735_ _3599_ _3736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6726_ _2240_ _2257_ _2837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4987_ _1072_ _1102_ _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6657_ _2680_ _2686_ _2769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6588_ _2700_ _2701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_116_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5608_ _1738_ _1740_ _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9108__CLK net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5539_ _1675_ _1676_ _1677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_8327_ _4096_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8258_ _4059_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9258__CLK net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7209_ _3262_ _3263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_6_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8189_ ci_adder.output_val_internal\[29\] ci_adder.output_val_internal\[21\] ci_adder.output_val_internal\[13\]
+ ci_adder.output_val_internal\[5\] _3964_ _3961_ _4016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_70_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5409__A1 _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4396__B2 internal_ih.byte0\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8288__I _4070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8685__I1 ci_adder.output_memory\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7637__A2 _3619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8775__CLK net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5890_ _2013_ _2014_ _2015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4910_ _0993_ _1063_ _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4841_ _0804_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_74_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7948__I0 _3718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6271__I _2388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4772_ _0898_ _0911_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7560_ _3552_ _3553_ _3554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4387__B2 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6511_ _2622_ _2624_ _2625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6128__A2 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8399__S _4122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7491_ _3496_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_31_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6442_ _2533_ _2556_ _2557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9230_ _0124_ net86 ci_adder.uut_simple_neuron.titan_id_5\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9161_ _0161_ net86 ci_adder.uut_simple_neuron.titan_id_3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6373_ _1950_ _1965_ _2489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8112_ _3804_ _3947_ _3950_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5639__A1 _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5324_ _1430_ _1457_ _1466_ _1467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9092_ _0545_ net34 ci_adder.output_val_internal\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5255_ _1263_ _1340_ _1399_ _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_11_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8043_ _3914_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5186_ _1298_ _1322_ _1331_ _1332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4862__A2 _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6064__A1 _2126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8945_ _0009_ net8 ci_adder.address_i\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8876_ _0423_ net63 ci_adder.output_memory\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7827_ _3778_ _3779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_104_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7564__A1 ci_adder.uut_simple_neuron.x0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4378__B2 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7758_ ci_adder.value_i\[21\] _3629_ _3722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6709_ _2818_ _2819_ _2820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7689_ _3487_ _3656_ _3664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8102__S _3825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9080__CLK net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8292__A2 _4071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4369__A1 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5869__A1 _1958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9054__D ci_adder.input_memory\[1\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8658__I1 ci_adder.output_memory\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8283__A2 _4071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5040_ _1157_ _1189_ _1190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7650__I _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6991_ ci_adder.uut_simple_neuron.titan_id_4\[18\] ci_adder.uut_simple_neuron.titan_id_3\[18\]
+ _3082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5942_ _2011_ _2022_ _2065_ _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_88_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7794__A1 _3632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8730_ net2 net43 spi_interface_cvonk.SS_r\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5873_ ci_adder.uut_simple_neuron.x3\[13\] ci_adder.uut_simple_neuron.x3\[14\] _1998_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_8661_ _4329_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8189__I3 ci_adder.output_val_internal\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4824_ _0956_ _0977_ _0979_ _0932_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8592_ ci_adder.uut_simple_neuron.x0\[26\] ci_adder.input_memory\[1\]\[26\] ci_adder.uut_simple_neuron.x2\[26\]
+ ci_adder.uut_simple_neuron.x3\[26\] _4252_ _4253_ _4285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7612_ _0688_ _3596_ _0684_ _3597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4755_ _0896_ _0912_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7543_ ci_adder.uut_simple_neuron.x0\[19\] _3539_ _3540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_43_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4686_ _0833_ _0838_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_9213_ _0079_ net38 ci_adder.uut_simple_neuron.titan_id_2\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7474_ _3481_ _3482_ _3483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6521__A2 _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6425_ _2471_ _2539_ _2540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_70_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9144_ _0236_ net91 ci_adder.uut_simple_neuron.titan_id_4\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6356_ _2365_ _2471_ _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5307_ _1445_ _1448_ _1450_ _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9075_ _0528_ net55 ci_adder.output_val_internal\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6287_ _1915_ _2404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8940__CLK net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8026_ _3905_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5238_ _1369_ _1383_ _1384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5169_ _1312_ _1315_ _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_8928_ _0001_ net10 ci_adder.address_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7936__S _3855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8859_ _0406_ net45 internal_ih.spi_tx_byte_o\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4771__A1 _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6028__A1 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8813__CLK net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4540_ ci_adder.uut_simple_neuron.x2\[0\] _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_53_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8963__CLK net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4471_ internal_ih.byte1\[4\] _0659_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6210_ _2118_ _2164_ _2329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7190_ _3245_ _3246_ _3247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4365__I1 internal_ih.byte3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6141_ _2242_ _2260_ _2261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9319__CLK net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6072_ _2141_ _2147_ _2193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5023_ _1134_ _1137_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4817__A2 ci_adder.uut_simple_neuron.x2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6019__A1 _1960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7767__A1 _3617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6974_ _3067_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5925_ ci_adder.uut_simple_neuron.x3\[12\] _1998_ _2048_ _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_88_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8713_ _0268_ net73 ci_adder.uut_simple_neuron.x3\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5856_ _1975_ _1977_ _1981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_101_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8644_ _4320_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _0960_ _0961_ _0962_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5787_ _1878_ _1880_ _1914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8582__I3 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8575_ _4257_ _4268_ _4270_ _4271_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4738_ _0875_ _0876_ _0895_ _0854_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_7526_ _3517_ _3522_ _3526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4669_ _0793_ _0828_ _0829_ _0715_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7457_ _3464_ _3467_ _3468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6408_ _2458_ _2521_ _2522_ _2523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_101_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9127_ ci_adder.uut_simple_neuron.x3\[0\] net86 ci_adder.uut_simple_neuron.titan_id_4\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7388_ _3407_ _3409_ _3410_ _3411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_112_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6339_ _1700_ _1702_ _2455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_112_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9058_ ci_adder.input_memory\[1\]\[26\] net28 ci_adder.uut_simple_neuron.titan_id_1\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4808__A2 _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8009_ _3896_ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6430__A1 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8836__CLK net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4441__B1 _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8986__CLK net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6249__A1 _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6544__I _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8410__A2 _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6421__A1 _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5710_ _1808_ _1811_ _1838_ _1839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6690_ _2754_ _2764_ _2800_ _2801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5641_ _1702_ _1755_ _1771_ _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__7772__I1 _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7921__A1 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5572_ _1696_ _1706_ _1707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4735__A1 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8360_ _4114_ _4109_ _4115_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7311_ _3346_ _3347_ _3348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8291_ _3452_ _4072_ _4078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4523_ ci_adder.address_i\[5\] ci_adder.address_i\[4\] ci_adder.address_i\[3\] _0693_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__8477__A2 _4170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9141__CLK net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7242_ ci_adder.uut_simple_neuron.titan_id_2\[28\] ci_adder.uut_simple_neuron.titan_id_5\[28\]
+ _3291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4454_ internal_ih.byte0\[4\] _0648_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5160__A1 _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7173_ _3231_ _3232_ _3233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8709__CLK net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4385_ _0614_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6124_ _2205_ _2208_ _2243_ _2244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6055_ _2173_ _2175_ _2176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9291__CLK net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5006_ _0831_ _0939_ _1082_ _1156_ _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__8859__CLK net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6957_ ci_adder.uut_simple_neuron.titan_id_4\[13\] ci_adder.uut_simple_neuron.titan_id_3\[13\]
+ _3053_ _3054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_49_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5908_ _2030_ _2031_ _1725_ _2032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6888_ _2949_ _2993_ _2996_ _2997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_62_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5839_ _1752_ _1964_ _1965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6715__A2 _2825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8627_ _0684_ _0687_ _0701_ _4311_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_36_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8558_ _4161_ _4257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_72_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7509_ _3510_ _3511_ _3512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8489_ ci_adder.output_memory\[8\] _4163_ _4200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5151__A1 _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9014__CLK net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4965__A1 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8156__A1 ci_adder.stream_o\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8546__I3 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5390__A1 _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7860_ internal_ih.spi_rx_byte_i\[2\] _3804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6811_ _2919_ _2920_ _2921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7198__A2 ci_adder.uut_simple_neuron.titan_id_5\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8490__S1 _4167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7791_ _3562_ _3730_ _3749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6742_ _2850_ _2852_ _2853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6673_ _2720_ _2781_ _2784_ _2785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_116_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5624_ _1702_ _1755_ _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_61_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8412_ _3733_ ci_adder.input_memory\[1\]\[23\] _4139_ _4144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8343_ _4104_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5555_ _1679_ ci_adder.uut_simple_neuron.x3\[3\] _1691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_124_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5486_ _1620_ _1625_ _1626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7122__A2 ci_adder.uut_simple_neuron.titan_id_5\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4506_ internal_ih.byte3\[5\] _0670_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8274_ _4067_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5133__A1 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4437_ internal_ih.byte6\[4\] _0635_ _0619_ internal_ih.byte2\[4\] _0644_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7225_ _3276_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7156_ ci_adder.uut_simple_neuron.titan_id_2\[15\] ci_adder.uut_simple_neuron.titan_id_5\[15\]
+ _3218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6107_ _1792_ _1810_ _2227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4368_ _0602_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_7087_ ci_adder.uut_simple_neuron.titan_id_2\[4\] ci_adder.uut_simple_neuron.titan_id_5\[4\]
+ _3160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6038_ _2156_ _2159_ _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__9037__CLK net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7189__A2 ci_adder.uut_simple_neuron.titan_id_5\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7989_ _3825_ _3886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9187__CLK net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7736__I1 ci_adder.uut_simple_neuron.x3\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7113__A2 ci_adder.uut_simple_neuron.titan_id_5\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6872__A1 _2974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8613__A2 _4301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6624__A1 ci_adder.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7975__I1 internal_ih.spi_rx_byte_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8015__S _3897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5340_ _0711_ _1448_ _1483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5271_ _1389_ _1415_ _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_23_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7010_ ci_adder.uut_simple_neuron.titan_id_4\[22\] ci_adder.uut_simple_neuron.titan_id_3\[22\]
+ _3097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6863__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8604__A2 _4161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8455__I2 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8961_ _0444_ net61 ci_adder.uut_simple_neuron.x0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_78_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7912_ _3840_ _3846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8892_ _0439_ net32 ci_adder.output_memory\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7843_ _3770_ _3791_ _3792_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout44_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4986_ _1134_ _1137_ _1138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4929__A1 _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7966__I1 ci_adder.uut_simple_neuron.x2\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7774_ ci_adder.uut_simple_neuron.x0\[24\] _3556_ _3726_ _3735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6725_ _2834_ _2835_ _2836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6656_ _2683_ _2685_ _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8540__A1 ci_adder.output_memory\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ _2648_ _2650_ _2699_ _2700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_104_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5607_ _1718_ _1739_ _1740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5538_ ci_adder.uut_simple_neuron.x3\[1\] _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8326_ _3723_ ci_adder.uut_simple_neuron.x0\[21\] _4091_ _4096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8257_ ci_adder.uut_simple_neuron.titan_id_6\[22\] _4059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5469_ _1573_ _1574_ _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7208_ ci_adder.uut_simple_neuron.titan_id_2\[23\] ci_adder.uut_simple_neuron.titan_id_5\[23\]
+ ci_adder.uut_simple_neuron.titan_id_2\[22\] ci_adder.uut_simple_neuron.titan_id_5\[22\]
+ _3262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_100_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8188_ _3963_ ci_adder.stream_o\[5\] ci_adder.stream_o\[21\] _3965_ _4014_ _4015_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_70_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7139_ ci_adder.uut_simple_neuron.titan_id_2\[12\] ci_adder.uut_simple_neuron.titan_id_5\[12\]
+ _3205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_6_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4396__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7709__I1 ci_adder.uut_simple_neuron.x3\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5345__A1 _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5648__A2 _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4840_ _0994_ _0983_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_117_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6510_ _1756_ _2623_ _2624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_99_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5584__A1 _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4771_ _0899_ _0874_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_56_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4387__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7490_ _3487_ _3493_ _3495_ _3496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_31_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6441_ _2551_ _2555_ _2556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6372_ _2483_ _2487_ _2488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9160_ _0160_ net86 ci_adder.uut_simple_neuron.titan_id_3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5323_ _1433_ _1456_ _1466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8111_ internal_ih.current_instruction\[2\] _3947_ _3950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9091_ _0544_ net34 ci_adder.output_val_internal\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5254_ _1221_ _1398_ _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_8042_ internal_ih.byte4\[1\] internal_ih.byte3\[1\] _3908_ _3914_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5185_ _1301_ _1321_ _1331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__9250__D _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8589__A1 ci_adder.output_val_internal\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8944_ _0008_ net8 ci_adder.address_i\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8875_ _0422_ net67 ci_adder.output_memory\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7826_ spi_interface_cvonk.SCLK_r\[2\] _3771_ _3773_ _3778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_47_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4969_ _0808_ _1083_ _1120_ _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4378__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7757_ _3539_ ci_adder.uut_simple_neuron.x0\[21\] _3715_ _3721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_117_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6708_ _2424_ _2659_ _2819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7688_ ci_adder.uut_simple_neuron.x0\[10\] _3657_ _3663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_116_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6639_ _2204_ _2750_ _2751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_59_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9225__CLK net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5878__A2 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8309_ _3680_ _3502_ _4076_ _4087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9289_ _0000_ net22 ci_adder.stream_enabled vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_83_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5566__A1 ci_adder.uut_simple_neuron.x3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8504__A1 ci_adder.output_memory\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5318__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5869__A2 _1960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6818__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8742__CLK net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6990_ _3065_ _3066_ _3080_ _3081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5941_ _2025_ _2064_ _2065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7794__A2 _3751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5872_ ci_adder.uut_simple_neuron.x3\[11\] _1959_ _1996_ _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_47_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8660_ ci_adder.stream_o\[15\] ci_adder.output_memory\[15\] _4323_ _4329_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4823_ _0978_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_16_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7611_ ci_adder.instruction_i\[2\] _3595_ _3596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_28_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8591_ ci_adder.output_memory\[26\] _4258_ _4284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4754_ _0898_ _0902_ _0911_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7542_ ci_adder.uut_simple_neuron.x0\[20\] _3539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_71_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7473_ _3480_ _3475_ _3478_ _3482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4685_ _0740_ _0789_ _0844_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_9212_ _0078_ net36 ci_adder.uut_simple_neuron.titan_id_2\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6424_ _2474_ _2538_ _2539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_70_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9143_ _0235_ net91 ci_adder.uut_simple_neuron.titan_id_4\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6355_ ci_adder.uut_simple_neuron.x3\[22\] _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6286_ _1694_ _2401_ _2402_ _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5306_ _0711_ _1449_ _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9074_ _0527_ net54 ci_adder.output_val_internal\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5237_ _1374_ _1376_ _1382_ _1383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7482__A1 _3479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8025_ internal_ih.byte3\[1\] internal_ih.byte2\[1\] _3897_ _3905_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ ci_adder.uut_simple_neuron.x2\[23\] _1267_ _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_3_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5099_ _1245_ _1247_ _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8927_ _0057_ net6 ci_adder.value_i\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8858_ _0405_ net44 internal_ih.spi_tx_byte_o\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8789_ _0336_ net41 internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7809_ ci_adder.uut_simple_neuron.x0\[30\] _3585_ _3754_ _3764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8113__S _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_117_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8765__CLK net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_58_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5787__A1 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8025__I0 internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7528__A2 _3524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_13_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8023__S _3897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4470_ _0661_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6140_ _2244_ _2259_ _2260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_96_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6071_ _1801_ _2191_ _2192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8693__S _3601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5022_ _1146_ _1172_ _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8492__I _4161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7767__A2 _3728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6973_ _3065_ _3066_ _3067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9070__CLK net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5924_ ci_adder.uut_simple_neuron.x3\[13\] ci_adder.uut_simple_neuron.x3\[14\] _2048_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_88_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8712_ _0267_ net73 ci_adder.uut_simple_neuron.x3\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__7519__A2 ci_adder.uut_simple_neuron.x0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4450__A1 internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5855_ _1980_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8643_ ci_adder.stream_o\[7\] ci_adder.output_memory\[7\] _4312_ _4320_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4806_ _0936_ _0907_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5786_ _1883_ _1887_ _1912_ _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_29_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8574_ ci_adder.output_val_internal\[22\] _4249_ _4271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5950__A1 _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4737_ _0712_ _0894_ _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7772__S _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7525_ ci_adder.uut_simple_neuron.x0\[15\] ci_adder.uut_simple_neuron.x0\[16\] _3525_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4668_ _0794_ _0817_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7456_ _3465_ _3466_ _3467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6407_ _2460_ _2499_ _2522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4599_ _0740_ _0762_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7387_ ci_adder.uut_simple_neuron.titan_id_1\[24\] ci_adder.uut_simple_neuron.titan_id_0\[24\]
+ _3410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9126_ _0192_ net26 ci_adder.uut_simple_neuron.titan_id_0\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6338_ _2452_ _2453_ _2454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_112_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7455__A1 ci_adder.uut_simple_neuron.x0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6269_ _2384_ _2386_ _2387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9057_ ci_adder.input_memory\[1\]\[25\] net28 ci_adder.uut_simple_neuron.titan_id_1\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8008_ internal_ih.byte2\[1\] internal_ih.byte1\[1\] _3886_ _3896_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_67_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7758__A2 _3629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4441__B2 internal_ih.byte2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4371__S _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8351__B _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6497__A2 _2364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7694__A1 _3617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9093__CLK net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6421__A2 _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8930__CLK net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5640_ _1752_ _1754_ _1771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7921__A2 _3846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5571_ _1699_ _1705_ _1706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7310_ ci_adder.uut_simple_neuron.titan_id_1\[11\] ci_adder.uut_simple_neuron.titan_id_0\[11\]
+ _3347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4522_ ci_adder.address_i\[17\] ci_adder.address_i\[16\] ci_adder.address_i\[15\]
+ ci_adder.address_i\[14\] _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_13_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8290_ _3454_ _4071_ _4077_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7241_ ci_adder.uut_simple_neuron.titan_id_2\[28\] ci_adder.uut_simple_neuron.titan_id_5\[28\]
+ _3290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7685__A1 _3619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4453_ _0652_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_84_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7172_ ci_adder.uut_simple_neuron.titan_id_2\[18\] ci_adder.uut_simple_neuron.titan_id_5\[18\]
+ _3232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4384_ internal_ih.byte7\[5\] _0603_ _0613_ net14 _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6123_ _2197_ _2204_ _2243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8485__I0 _3470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6054_ _2174_ _2129_ _2175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout74_I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6660__A2 _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5005_ _0831_ _0939_ _1112_ _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__8155__C _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_93_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6956_ _3049_ _3050_ _3052_ _3053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_88_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5907_ _1709_ _1990_ _2031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__B2 internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6887_ _2994_ _2938_ _2995_ _2937_ _2996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_118_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5838_ _1754_ _1843_ _1964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_76_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8626_ _0684_ _0687_ ci_adder.interrupt_enabled _4311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5769_ _1896_ _1856_ _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5923__A1 _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8557_ _4211_ _4251_ _4255_ _4256_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7508_ ci_adder.uut_simple_neuron.x0\[11\] _3502_ ci_adder.uut_simple_neuron.x0\[12\]
+ _3511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_16_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7676__A1 _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8488_ _4162_ _4196_ _4198_ _4199_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_102_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7439_ ci_adder.uut_simple_neuron.x0\[4\] _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_32_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9109_ _0174_ net60 ci_adder.uut_simple_neuron.titan_id_0\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8803__CLK net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8953__CLK net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6167__A1 _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9309__CLK net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8301__S _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7667__A1 ci_adder.uut_simple_neuron.x3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6810_ _0162_ _2853_ _2920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4405__A1 internal_ih.byte4\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4405__B2 internal_ih.byte0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7790_ ci_adder.value_i\[27\] _3629_ _3748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6741_ _1836_ _2851_ _2852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6672_ _2648_ _2782_ _2783_ _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5623_ _1752_ _1754_ _1755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_8411_ _3728_ _4117_ _4143_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8342_ _3762_ ci_adder.uut_simple_neuron.x0\[29\] _4070_ _4104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5554_ _1675_ _1688_ _1689_ _1690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_6_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7658__A1 _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5485_ _1481_ _1624_ _1625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__9253__D _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4505_ _0679_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8273_ ci_adder.uut_simple_neuron.titan_id_6\[30\] _4067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7224_ _3274_ _3275_ _3276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4436_ _0643_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8826__CLK net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8010__I _3825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7155_ _3217_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4367_ internal_ih.current_instruction\[1\] _0601_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6106_ _2185_ _2211_ _2225_ _2226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7086_ _3159_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6037_ _2033_ _2157_ _2158_ _2159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8976__CLK net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8386__A2 _4117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7988_ _3885_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6939_ ci_adder.uut_simple_neuron.titan_id_4\[10\] ci_adder.uut_simple_neuron.titan_id_3\[10\]
+ _3039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_49_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7897__A1 _3826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8609_ ci_adder.output_val_internal\[29\] _4161_ _4299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8449__I0 ci_adder.uut_simple_neuron.x0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8377__A2 _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9131__CLK net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6560__A1 _2249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5270_ _1392_ _1394_ _1414_ _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_120_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8455__I3 _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8960_ _0443_ net41 internal_ih.received_byte_count\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7911_ _3625_ _3841_ _3845_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8891_ _0438_ net32 ci_adder.output_memory\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8368__A2 _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7842_ internal_ih.spi_rx_byte_i\[3\] _3787_ _3792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4985_ _0996_ _1135_ _1136_ _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9248__D _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7773_ _3734_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout37_I net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6724_ _2197_ _2751_ _2835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6655_ _2694_ _2695_ _2767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_12_Left_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8540__A2 _4212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ _2689_ _2698_ _2699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6551__A1 _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5606_ _1716_ _1739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5537_ ci_adder.uut_simple_neuron.x3\[0\] _1675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_8325_ _4095_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8256_ _4058_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5468_ _1606_ _1607_ _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7207_ _3254_ _3259_ _3261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5399_ _1518_ _1540_ _1541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4419_ _0634_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8187_ _3966_ _4013_ _4014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7138_ _3200_ _3202_ _3203_ _3204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_6_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7069_ _3144_ _3145_ _3146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9154__CLK net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9158__D ci_adder.uut_simple_neuron.x2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5345__A2 ci_adder.uut_simple_neuron.x2\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8295__A1 _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7098__A2 ci_adder.uut_simple_neuron.titan_id_5\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5648__A3 _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6845__A2 ci_adder.uut_simple_neuron.x3\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8598__A2 _4289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4608__A1 _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7929__I _3840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5033__A1 _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6781__A1 ci_adder.uut_simple_neuron.x3\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4770_ _0834_ _0926_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_67_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6440_ _2047_ _2554_ _2555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6371_ _1995_ _2486_ _2487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9027__CLK net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5322_ _1465_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8110_ _3949_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9090_ _0543_ net34 ci_adder.output_val_internal\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5253_ _1233_ ci_adder.uut_simple_neuron.x2\[22\] ci_adder.uut_simple_neuron.x2\[23\]
+ _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_11_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8041_ _3913_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9177__CLK net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5184_ _0994_ _1324_ _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5272__A1 _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8943_ _0007_ net8 ci_adder.address_i\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8874_ _0421_ net67 ci_adder.output_memory\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7825_ _3775_ _3777_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_50_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7775__S _3599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4968_ _1016_ _1057_ _1095_ _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_62_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7756_ _3539_ _3715_ ci_adder.uut_simple_neuron.x0\[21\] _3720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6707_ _2468_ _2599_ _2818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4899_ _0811_ _1052_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7687_ _3662_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6524__A1 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6638_ _2300_ _2748_ _2749_ _2750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_6_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8513__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4386__I0 internal_ih.byte4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6569_ _2094_ _2613_ _2682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8308_ _4086_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9288_ _0550_ net23 ci_adder.interrupt_enabled vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8239_ ci_adder.uut_simple_neuron.titan_id_6\[13\] _4050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7252__A2 ci_adder.uut_simple_neuron.titan_id_5\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4374__S _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_83_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6763__A1 _2797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5566__A2 ci_adder.uut_simple_neuron.x3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6515__A1 _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8504__A2 _4212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4377__I0 internal_ih.byte4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5940_ _2026_ _2063_ _2064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_36_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5871_ ci_adder.uut_simple_neuron.x3\[12\] ci_adder.uut_simple_neuron.x3\[13\] _1996_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_87_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5006__A1 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7610_ _0685_ _0686_ _3595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4822_ _0714_ _0976_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_8_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_16_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8590_ _4257_ _4280_ _4282_ _4283_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4753_ _0852_ _0910_ _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_71_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7541_ _3538_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7472_ _3475_ _3478_ _3480_ _3481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4684_ _0785_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_9211_ _0076_ net74 ci_adder.uut_simple_neuron.titan_id_2\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6423_ ci_adder.uut_simple_neuron.x3\[24\] _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_43_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6354_ _2252_ _2425_ _2469_ _2470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9142_ _0234_ net88 ci_adder.uut_simple_neuron.titan_id_4\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6285_ _1909_ _2348_ _2402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5305_ _1404_ _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_9073_ _0526_ net57 ci_adder.output_val_internal\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5236_ _1326_ _1378_ _1380_ _1381_ _1382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7482__A2 ci_adder.uut_simple_neuron.x0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8024_ _3904_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ _1310_ _1311_ _1313_ _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5098_ _1198_ _1208_ _1246_ _1247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5245__A1 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8926_ _0056_ net6 ci_adder.value_i\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8857_ _0404_ net46 internal_ih.spi_tx_byte_o\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6745__A1 _2844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8788_ _0335_ net42 internal_ih.byte0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7808_ _3763_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7739_ _3531_ _3695_ _3706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_104_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_113_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5787__A2 _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6984__A1 ci_adder.uut_simple_neuron.titan_id_4\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8025__I1 internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5539__A2 _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8489__A1 ci_adder.output_memory\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6070_ _1807_ _2190_ _2191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5475__A1 _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5021_ _0993_ _1171_ _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_49_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6972_ ci_adder.uut_simple_neuron.titan_id_4\[16\] ci_adder.uut_simple_neuron.titan_id_3\[16\]
+ _3066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6975__A1 ci_adder.uut_simple_neuron.titan_id_4\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8711_ _0266_ net74 ci_adder.uut_simple_neuron.x3\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5923_ _1880_ _2000_ _2046_ _2047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_76_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5854_ _1941_ _1942_ _1979_ _1980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__6727__A1 _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8567__I2 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8642_ _4319_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4805_ _0936_ _0907_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8573_ _4260_ _4269_ _4270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5785_ _1876_ _1882_ _1912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4541__I _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7524_ ci_adder.uut_simple_neuron.x0\[17\] _3524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_16_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5950__A2 _2072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4736_ ci_adder.uut_simple_neuron.x2\[9\] ci_adder.uut_simple_neuron.x2\[10\] ci_adder.uut_simple_neuron.x2\[11\]
+ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4667_ _0802_ _0817_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7455_ ci_adder.uut_simple_neuron.x0\[3\] _3459_ _3452_ _3466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_31_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6406_ _2460_ _2499_ _2521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7386_ ci_adder.uut_simple_neuron.titan_id_1\[24\] ci_adder.uut_simple_neuron.titan_id_0\[24\]
+ _3409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6337_ _2403_ _2409_ _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4598_ _0749_ _0752_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9125_ _0191_ net25 ci_adder.uut_simple_neuron.titan_id_0\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6268_ _2318_ _2385_ _2386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9056_ ci_adder.input_memory\[1\]\[24\] net29 ci_adder.uut_simple_neuron.titan_id_1\[26\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7455__A2 _3459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6199_ _2314_ _2317_ _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5219_ _0996_ _1364_ _1365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8007_ _3895_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8909_ _0037_ net12 ci_adder.value_i\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8732__CLK net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4451__I _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8882__CLK net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8034__S _3908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5570_ _1704_ _1705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4521_ ci_adder.address_i\[13\] ci_adder.address_i\[12\] ci_adder.address_i\[11\]
+ ci_adder.address_i\[10\] _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_13_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4452_ internal_ih.byte0\[3\] _0648_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7240_ _3289_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4743__I0 _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7171_ ci_adder.uut_simple_neuron.titan_id_2\[17\] ci_adder.uut_simple_neuron.titan_id_5\[17\]
+ _3220_ _3228_ _3230_ _3231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4383_ internal_ih.byte4\[5\] internal_ih.byte3\[5\] _0599_ _0613_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6122_ _1841_ _2241_ _2242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7437__A2 ci_adder.uut_simple_neuron.x0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6053_ _1723_ _1757_ _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5004_ _1122_ _1129_ _1154_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4671__A2 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout67_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7996__I0 internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6955_ ci_adder.uut_simple_neuron.titan_id_4\[12\] ci_adder.uut_simple_neuron.titan_id_3\[12\]
+ _3052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_89_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5906_ _1715_ _1989_ _2030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5620__A1 ci_adder.uut_simple_neuron.x3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__A2 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6886_ _2870_ _2867_ _2995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_62_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7748__I0 _3713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8625_ _4310_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5837_ _1956_ _1962_ _1963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_57_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5768_ _1828_ _1816_ _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_106_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8556_ ci_adder.output_val_internal\[19\] _4249_ _4256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4719_ _0718_ _0852_ _0856_ _0849_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_72_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7507_ ci_adder.uut_simple_neuron.x0\[12\] _3502_ _3498_ _3499_ _3497_ _3510_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_8487_ ci_adder.output_val_internal\[7\] _4170_ _4199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5699_ _1781_ _1784_ _1828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7438_ _3451_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7369_ ci_adder.uut_simple_neuron.titan_id_1\[21\] ci_adder.uut_simple_neuron.titan_id_0\[21\]
+ _3396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9108_ _0173_ net58 ci_adder.uut_simple_neuron.titan_id_0\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9039_ ci_adder.input_memory\[1\]\[7\] net65 ci_adder.uut_simple_neuron.titan_id_1\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7958__S _3840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7987__I0 internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5611__A1 _1735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__A1 _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7667__A2 _3617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9060__CLK net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8616__A1 ci_adder.output_memory\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8029__S _3897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8778__CLK net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8475__S0 _4166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6740_ _1841_ _1851_ _2851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4405__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6671_ _2650_ _2699_ _2783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5622_ ci_adder.uut_simple_neuron.x3\[5\] _1753_ _1754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_8410_ ci_adder.input_memory\[1\]\[22\] _4118_ _4143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5553_ _1676_ _1679_ _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8341_ _4103_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4504_ internal_ih.byte3\[4\] _0670_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_26_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5484_ _1479_ _1623_ _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8272_ _4066_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7658__A2 _3459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7223_ ci_adder.uut_simple_neuron.titan_id_2\[26\] ci_adder.uut_simple_neuron.titan_id_5\[26\]
+ _3275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4435_ internal_ih.byte6\[3\] _0635_ _0632_ internal_ih.byte2\[3\] _0643_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7154_ ci_adder.uut_simple_neuron.titan_id_2\[15\] ci_adder.uut_simple_neuron.titan_id_5\[15\]
+ _3216_ _3217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4366_ _0597_ _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6105_ _2188_ _2210_ _2225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7085_ _3157_ _3158_ _3159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6036_ _2076_ _2110_ _2158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_83_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7987_ internal_ih.byte0\[7\] internal_ih.spi_rx_byte_i\[7\] _3877_ _3885_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_1_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6938_ ci_adder.uut_simple_neuron.titan_id_4\[9\] ci_adder.uut_simple_neuron.titan_id_3\[9\]
+ _3035_ _3036_ _3038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_120_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6869_ _2292_ _2307_ _2978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4930__S _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8608_ _4260_ _4297_ _4298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9083__CLK net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8539_ _4211_ _4238_ _4240_ _4241_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_103_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4580__A1 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4377__S _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6085__A1 _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8920__CLK net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__A1 ci_adder.uut_simple_neuron.x3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7487__I ci_adder.uut_simple_neuron.x0\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4399__B2 internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6076__A1 _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7910_ _0724_ _3842_ _3845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8890_ _0437_ net32 ci_adder.output_memory\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7841_ internal_ih.spi_tx_byte_o\[2\] _3779_ _3784_ internal_ih.spi_rx_byte_i\[2\]
+ _3791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4984_ _1075_ _1100_ _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7772_ _3733_ _2474_ _3692_ _3734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6723_ _2204_ _2750_ _2834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6654_ _2725_ _2765_ _2766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_74_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5605_ _1722_ _1735_ _1737_ _1738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_73_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6585_ _2690_ _2697_ _2698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5536_ _1674_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4562__A1 _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8324_ _3718_ _3539_ _4091_ _4095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8679__I1 ci_adder.output_memory\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5467_ _1482_ _1576_ _1607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8943__CLK net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8255_ ci_adder.uut_simple_neuron.titan_id_6\[21\] _4058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4418_ internal_ih.byte5\[3\] _0623_ _0632_ internal_ih.byte1\[3\] _0634_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7206_ _3260_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5398_ _1437_ _1539_ _1540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8186_ _3962_ ci_adder.stream_o\[13\] _4013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_70_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7137_ ci_adder.uut_simple_neuron.titan_id_2\[11\] ci_adder.uut_simple_neuron.titan_id_5\[11\]
+ _3203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4349_ _0583_ internal_ih.received_byte_count\[2\] internal_ih.expected_byte_count\[3\]
+ _0584_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7068_ ci_adder.uut_simple_neuron.titan_id_2\[1\] ci_adder.uut_simple_neuron.titan_id_5\[1\]
+ _3145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6019_ _1960_ _2101_ _2140_ _2141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_68_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8295__A2 _4072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7703__C _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6058__A1 _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4608__A2 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8307__S _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8816__CLK net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6781__A2 ci_adder.uut_simple_neuron.x3\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8042__S _3908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8602__S0 _4252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8966__CLK net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _2001_ _2485_ _2486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5321_ _1463_ _1464_ _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8040_ internal_ih.byte4\[0\] internal_ih.byte3\[0\] _3908_ _3913_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8286__A2 _4072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5252_ _1395_ _1358_ _1396_ _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5183_ _1296_ _1323_ _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8942_ _0006_ net8 ci_adder.address_i\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8873_ _0420_ net63 ci_adder.output_memory\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4544__I _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7824_ net5 _3776_ _3777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4967_ _0808_ _1083_ _1080_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7755_ _2467_ _3612_ _3719_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6706_ _2808_ _2816_ _2817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4898_ _1049_ _1051_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7686_ _3661_ ci_adder.uut_simple_neuron.x3\[9\] _3632_ _3662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6637_ _2302_ _2545_ _2749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7721__A1 _3619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_119_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6568_ _2102_ _2612_ _2681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5519_ _1654_ _1657_ _1658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8307_ _3677_ ci_adder.uut_simple_neuron.x0\[12\] _4076_ _4086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6499_ _2102_ _2612_ _2613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6288__A1 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9287_ _0549_ net32 ci_adder.normalised_stream_write_address\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8238_ _4049_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8169_ _3966_ _3997_ _3998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8839__CLK net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7966__S _3840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6212__A1 _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7960__A1 _3746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8989__CLK net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4774__A1 _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6515__A2 _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6844__I ci_adder.uut_simple_neuron.x3\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5870_ _1845_ _1961_ _1994_ _1995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_87_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4821_ _0976_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5006__A2 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4765__A1 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4752_ _0814_ _0909_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7540_ _3536_ _3537_ _3538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_126_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4683_ _0843_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7471_ _3470_ _3479_ _3480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9144__CLK net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6422_ _2365_ _2475_ _2536_ _2537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_9210_ _0075_ net74 ci_adder.uut_simple_neuron.titan_id_2\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9141_ _0233_ net88 ci_adder.uut_simple_neuron.titan_id_4\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6353_ _2422_ _2468_ _2469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_12_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6284_ _1909_ _2348_ _2401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5304_ _1442_ _1446_ _1447_ _1448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_59_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9072_ _0525_ net56 ci_adder.output_val_internal\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5235_ _1293_ _1377_ _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8023_ internal_ih.byte3\[0\] internal_ih.byte2\[0\] _3897_ _3904_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5166_ _1233_ _1312_ _1313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5097_ _1194_ _1197_ _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8925_ _0054_ net6 ci_adder.value_i\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8856_ _0403_ net42 internal_ih.spi_tx_byte_o\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5999_ _2085_ _2108_ _2121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8787_ _0334_ net42 internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7807_ _3762_ ci_adder.uut_simple_neuron.x3\[29\] _3611_ _3763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7738_ ci_adder.value_i\[18\] _3629_ _3705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7669_ _3469_ _3470_ _3638_ _3647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_30_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6681__A1 _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9017__CLK net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4995__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9167__CLK net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4747__A1 ci_adder.uut_simple_neuron.x2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8320__S _4091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5172__A1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6672__A1 _2648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5020_ _1149_ _1170_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5475__A2 ci_adder.uut_simple_neuron.x2\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6424__A1 _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ _3061_ _3063_ _3064_ _3065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8710_ _0265_ net74 ci_adder.uut_simple_neuron.x3\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_49_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5922_ _1997_ _1999_ _2046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5853_ _1975_ _1978_ _1979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_76_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7924__A1 _3654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8567__I3 _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8641_ ci_adder.stream_o\[6\] ci_adder.output_memory\[6\] _4312_ _4319_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5784_ _1695_ _1910_ _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4804_ _0904_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_75_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8572_ ci_adder.uut_simple_neuron.x0\[22\] ci_adder.input_memory\[1\]\[22\] ci_adder.uut_simple_neuron.x2\[22\]
+ _2471_ _4252_ _4253_ _4269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_91_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4735_ _0811_ _0834_ _0852_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7523_ _3523_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout12_I internal_ih.got_all_data vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4666_ _0804_ _0819_ _0826_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7152__A2 ci_adder.uut_simple_neuron.titan_id_5\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7454_ _3452_ _3459_ _3453_ _3457_ _3465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6405_ _2519_ _2520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_101_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4597_ _0759_ _0760_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7385_ _3408_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6336_ _2406_ _2408_ _2452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4910__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9124_ _0189_ net27 ci_adder.uut_simple_neuron.titan_id_0\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9055_ ci_adder.input_memory\[1\]\[23\] net29 ci_adder.uut_simple_neuron.titan_id_1\[25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6267_ _2269_ _2268_ _2385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6198_ _2315_ _2264_ _2316_ _2317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5218_ _1332_ _1363_ _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8006_ internal_ih.byte2\[0\] internal_ih.byte1\[0\] _3886_ _3895_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5149_ _1251_ _1294_ _1295_ _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_67_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8908_ _0036_ net12 ci_adder.value_i\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7915__A1 ci_adder.uut_simple_neuron.x2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8839_ _0386_ net21 internal_ih.byte7\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6394__I _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4968__A1 _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8315__S _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7906__A1 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4520_ ci_adder.address_i\[21\] ci_adder.address_i\[20\] ci_adder.address_i\[19\]
+ ci_adder.address_i\[18\] _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__8050__S _3908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5145__A1 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4451_ _0651_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7170_ _3229_ _3230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6121_ _1847_ _2240_ _2241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4382_ _0612_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8485__I2 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6052_ _2125_ _2128_ _2173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_111_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5003_ _1123_ _1128_ _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6954_ _3051_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5905_ _1985_ _2027_ _2028_ _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6885_ _2792_ _2865_ _2994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_118_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7748__I1 _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8624_ _4167_ ci_adder.normalised_stream_write_address\[1\] _4308_ _4310_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5836_ _1845_ _1961_ _1962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_62_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5767_ _1866_ _1891_ _1894_ _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8555_ _4214_ _4254_ _4255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5698_ _1764_ _1819_ _1826_ _1816_ _1827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4718_ _0875_ _0876_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7506_ _3502_ _3508_ _3509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_17_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8486_ _4165_ _4197_ _4198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4649_ _0740_ _0790_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_0_71_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7437_ _3447_ ci_adder.uut_simple_neuron.x0\[3\] _3450_ _3451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_102_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7368_ _3391_ _3392_ _3394_ _3395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6319_ _2413_ _2435_ _2436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7299_ ci_adder.uut_simple_neuron.titan_id_1\[9\] ci_adder.uut_simple_neuron.titan_id_0\[9\]
+ _3337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9107_ _0172_ net58 ci_adder.uut_simple_neuron.titan_id_0\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9038_ ci_adder.input_memory\[1\]\[6\] net67 ci_adder.uut_simple_neuron.titan_id_1\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7833__B1 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7987__I1 internal_ih.spi_rx_byte_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_43_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5678__A2 _1807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8616__A2 _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8475__S1 _4167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6670_ _2650_ _2699_ _2782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5621_ ci_adder.uut_simple_neuron.x3\[6\] ci_adder.uut_simple_neuron.x3\[7\] _1753_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_45_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7683__I _3608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5552_ _1676_ _1679_ _1688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8340_ _3757_ ci_adder.uut_simple_neuron.x0\[28\] _4070_ _4103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5118__A1 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4503_ _0678_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8271_ ci_adder.uut_simple_neuron.titan_id_6\[29\] _4066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5483_ _1572_ _1621_ _1622_ _1623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7222_ _3267_ _3271_ _3273_ _3274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4434_ _0642_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7153_ _3212_ _3213_ _3215_ _3216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4365_ internal_ih.byte4\[0\] internal_ih.byte3\[0\] _0599_ _0600_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6104_ _2222_ _2223_ _2224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7084_ ci_adder.uut_simple_neuron.titan_id_2\[4\] ci_adder.uut_simple_neuron.titan_id_5\[4\]
+ _3158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6035_ _2076_ _2110_ _2157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8722__CLK net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7986_ _3884_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8182__C _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8872__CLK net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6937_ _3037_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6868_ _2975_ _2976_ _2977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5819_ _1943_ _1944_ _1945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5357__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8607_ ci_adder.uut_simple_neuron.x0\[29\] ci_adder.input_memory\[1\]\[29\] ci_adder.uut_simple_neuron.x2\[29\]
+ ci_adder.uut_simple_neuron.x3\[29\] _0698_ _0697_ _4297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_6799_ _2254_ _2825_ _2909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8538_ ci_adder.output_val_internal\[16\] _4203_ _4241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5109__A1 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4580__A2 _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8469_ ci_adder.output_memory\[4\] _4163_ _4184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8449__I2 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5596__A1 ci_adder.uut_simple_neuron.x3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4399__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8534__A1 _4211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_97_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4626__A3 ci_adder.uut_simple_neuron.x2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8895__CLK net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7840_ _3770_ _3789_ _3790_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8612__I2 ci_adder.uut_simple_neuron.x2\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4983_ _1075_ _1100_ _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7771_ _3619_ _3730_ _3731_ _3732_ _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_106_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6722_ _2831_ _2832_ _2833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8525__A1 ci_adder.output_memory\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6653_ _2754_ _2764_ _2765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5604_ _1678_ _1716_ _1736_ _1737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_74_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6584_ _2693_ _2696_ _2697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_26_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5535_ _1663_ _1671_ _1673_ _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_5_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8323_ _4094_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_124_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6839__A1 _2349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5466_ _1566_ _1567_ _1575_ _1606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8254_ _4057_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5511__A1 _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7205_ _3258_ _3259_ _3260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4417_ _0633_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5397_ _1521_ _1538_ _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8185_ _3979_ _4011_ _4012_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_70_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7136_ ci_adder.uut_simple_neuron.titan_id_2\[11\] ci_adder.uut_simple_neuron.titan_id_5\[11\]
+ _3202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_6_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4348_ internal_ih.received_byte_count\[3\] _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7067_ ci_adder.uut_simple_neuron.titan_id_2\[0\] ci_adder.uut_simple_neuron.titan_id_5\[0\]
+ _3144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6018_ _2097_ _2100_ _2140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_94_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5578__A1 ci_adder.uut_simple_neuron.x3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9050__CLK net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7969_ _3875_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5750__A1 ci_adder.uut_simple_neuron.x3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7699__S _3632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8055__I0 internal_ih.byte4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7558__A2 ci_adder.uut_simple_neuron.x0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8602__S1 _4253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5320_ _1418_ _1423_ _1419_ _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5251_ _0714_ _1316_ _1356_ _1396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_11_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ _1328_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_3_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8941_ _0005_ net7 ci_adder.address_i\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_108_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8046__I0 internal_ih.byte4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9073__CLK net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8872_ _0419_ net63 ci_adder.output_memory\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7823_ _3770_ _3772_ _3776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout42_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7754_ _3632_ _3718_ _3719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6705_ _2601_ _2815_ _2816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4966_ _1088_ _1097_ _1117_ _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_50_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4783__A2 _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4897_ _0909_ _0939_ _1050_ _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_62_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7685_ _3619_ _3657_ _3658_ _3660_ _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_46_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8910__CLK net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6636_ _2302_ _2545_ _2748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_119_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6567_ _2678_ _2679_ _2680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5518_ _1560_ _1655_ _1656_ _1657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8306_ _3493_ _4071_ _4085_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6498_ _2199_ _2549_ _2611_ _2612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9286_ _0548_ net22 ci_adder.normalised_stream_write_address\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5449_ _1513_ _1547_ _1590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8237_ ci_adder.uut_simple_neuron.titan_id_6\[12\] _4049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8168_ _3962_ ci_adder.stream_o\[11\] _3997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7119_ ci_adder.uut_simple_neuron.titan_id_2\[9\] ci_adder.uut_simple_neuron.titan_id_5\[9\]
+ _3188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8408__S _4139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8099_ _3943_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4471__A1 internal_ih.byte1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__A2 _2072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7960__A2 _3846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5971__A1 _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__A2 ci_adder.uut_simple_neuron.x2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7476__A1 _3470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8318__S _4091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4820_ _0874_ _0975_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8053__S _3919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4751_ _0908_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9095__D ci_adder.uut_simple_neuron.x0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4682_ _0824_ _0827_ _0842_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__8587__S0 _4252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7470_ ci_adder.uut_simple_neuron.x0\[8\] _3479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_43_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6421_ _2471_ _2474_ _2536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5714__A1 ci_adder.uut_simple_neuron.x3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9140_ _0232_ net89 ci_adder.uut_simple_neuron.titan_id_4\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6352_ _2467_ _2423_ _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6283_ _2351_ _2374_ _2399_ _2400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5303_ ci_adder.uut_simple_neuron.x2\[24\] ci_adder.uut_simple_neuron.x2\[25\] ci_adder.uut_simple_neuron.x2\[26\]
+ _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__7467__A1 _3459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9071_ _0524_ net56 ci_adder.output_val_internal\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5234_ _1288_ _1379_ _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8022_ _3903_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6690__A2 _2764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5165_ _1221_ _1268_ _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8511__S0 _4206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5096_ _1243_ _1244_ _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8924_ _0053_ net6 ci_adder.value_i\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8019__I0 internal_ih.byte2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6993__A3 _3083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8855_ _0402_ net41 internal_ih.instruction_received vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_93_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7806_ _3659_ _3759_ _3760_ _3761_ _3762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_5998_ _2079_ _2080_ _2081_ _2120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_93_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8786_ _0333_ net19 internal_ih.byte0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4949_ _0870_ _1101_ _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7737_ _3704_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7668_ _3612_ _3645_ _3646_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6619_ _2729_ _2730_ _2731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4508__A2 _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7599_ ci_adder.uut_simple_neuron.x0\[28\] ci_adder.uut_simple_neuron.x0\[29\] _3586_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9269_ _0133_ net82 ci_adder.uut_simple_neuron.titan_id_6\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_18_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8806__CLK net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8956__CLK net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7630__A1 ci_adder.uut_simple_neuron.x0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5944__A1 _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7697__A1 ci_adder.value_i\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5172__A2 _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6121__A1 _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8048__S _3908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6424__A2 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6970_ ci_adder.uut_simple_neuron.titan_id_4\[15\] ci_adder.uut_simple_neuron.titan_id_3\[15\]
+ _3064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_45_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _2002_ _2005_ _2044_ _2045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4435__B2 internal_ih.byte2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5852_ _1976_ _1977_ _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6188__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7924__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9111__CLK net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8640_ _4318_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5783_ _1907_ _1909_ _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4803_ _0900_ _0956_ _0958_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8571_ ci_adder.output_memory\[22\] _4258_ _4268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4734_ _0872_ _0879_ _0880_ _0882_ _0804_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_7522_ _3517_ _3522_ _3523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4665_ _0770_ _0825_ _0818_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_54_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7453_ _3459_ ci_adder.uut_simple_neuron.x0\[6\] _3464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6404_ _2452_ _2453_ _2457_ _2519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_116_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6360__A1 _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4596_ _0738_ _0755_ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7384_ ci_adder.uut_simple_neuron.titan_id_1\[24\] ci_adder.uut_simple_neuron.titan_id_0\[24\]
+ _3407_ _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_3_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8829__CLK net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6335_ _2398_ _2438_ _2450_ _2451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_101_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5155__B _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9123_ _0188_ net31 ci_adder.uut_simple_neuron.titan_id_0\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6112__A1 _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9054_ ci_adder.input_memory\[1\]\[22\] net29 ci_adder.uut_simple_neuron.titan_id_1\[24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6266_ _2321_ _2333_ _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8005_ _3894_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6197_ _2226_ _2263_ _2316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5217_ _1335_ _1362_ _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4674__A1 _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5148_ _1256_ _1278_ _1295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_63_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5079_ _1225_ _1227_ _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_67_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8907_ _0035_ net12 ci_adder.value_i\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6179__A1 _2100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8412__I0 _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8838_ _0385_ net15 internal_ih.byte6\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8769_ _0316_ net73 ci_adder.uut_simple_neuron.x2\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7915__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7679__A1 _3612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6103__A1 _2126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9134__CLK net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7906__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7455__B _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4450_ internal_ih.byte0\[2\] _0648_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4381_ internal_ih.byte7\[4\] _0603_ _0611_ net14 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_111_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6120_ _1917_ _2206_ _2239_ _2240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__8485__I3 ci_adder.uut_simple_neuron.x3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6051_ _2120_ _2170_ _2171_ _2172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_111_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7842__A1 internal_ih.spi_rx_byte_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5002_ _1084_ _1120_ _1152_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_95_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6953_ _3049_ _3050_ _3051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4959__A2 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5904_ _1987_ _2007_ _2028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6884_ _2962_ _2983_ _2992_ _2993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_88_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5835_ _1958_ _1960_ _1961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_64_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8623_ _4309_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_62_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5766_ _1793_ _1892_ _1893_ _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8554_ ci_adder.uut_simple_neuron.x0\[19\] ci_adder.input_memory\[1\]\[19\] ci_adder.uut_simple_neuron.x2\[19\]
+ _2250_ _4252_ _4253_ _4254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_44_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5697_ _1781_ _1784_ _1826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4717_ _0849_ _0852_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8485_ _3470_ ci_adder.input_memory\[1\]\[7\] _0787_ ci_adder.uut_simple_neuron.x3\[7\]
+ _4166_ _4167_ _4197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_7505_ ci_adder.uut_simple_neuron.x0\[14\] _3508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6333__A1 _1721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4648_ _0806_ _0808_ _0809_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7436_ ci_adder.uut_simple_neuron.x0\[2\] _3448_ _3450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9007__CLK net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4895__A1 _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4579_ _0739_ _0743_ _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9106_ _0171_ net65 ci_adder.uut_simple_neuron.titan_id_0\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7367_ ci_adder.uut_simple_neuron.titan_id_1\[20\] ci_adder.uut_simple_neuron.titan_id_0\[20\]
+ _3394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6318_ _2430_ _2434_ _2435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7298_ _3336_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6249_ _2250_ _2366_ _2367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4647__A1 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9037_ ci_adder.input_memory\[1\]\[5\] net66 ci_adder.uut_simple_neuron.titan_id_1\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7833__B2 internal_ih.spi_rx_byte_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9157__CLK net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8416__S _4139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6572__A1 _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6324__A1 _2391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6875__A2 _2931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8624__I0 _4167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8326__S _4091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5620_ ci_adder.uut_simple_neuron.x3\[4\] _1731_ _1751_ _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__8061__S _3919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5551_ _1679_ ci_adder.uut_simple_neuron.x3\[3\] _1687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_124_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8304__A2 _4072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4502_ internal_ih.byte3\[3\] _0670_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8270_ _4065_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5482_ ci_adder.uut_simple_neuron.x2\[27\] _1530_ _1569_ _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7221_ _3268_ _3273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4433_ internal_ih.byte6\[2\] _0635_ _0632_ internal_ih.byte2\[2\] _0642_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7152_ ci_adder.uut_simple_neuron.titan_id_2\[14\] ci_adder.uut_simple_neuron.titan_id_5\[14\]
+ _3215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4364_ _0598_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6103_ _2126_ _2184_ _2223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7083_ _3154_ _3156_ _3157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6034_ _2120_ _2122_ _2155_ _2156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__4629__A1 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout72_I net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7985_ internal_ih.byte0\[6\] internal_ih.spi_rx_byte_i\[6\] _3877_ _3884_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6936_ _3035_ _3036_ _3037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6867_ _2918_ _2933_ _2976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8543__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5818_ _1682_ _1910_ _1944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6798_ _2906_ _2907_ _2908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8606_ ci_adder.output_memory\[29\] _4258_ _4296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5749_ ci_adder.uut_simple_neuron.x3\[9\] ci_adder.uut_simple_neuron.x3\[10\] _1877_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_45_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8537_ _4214_ _4239_ _4240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_20_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4580__A3 ci_adder.uut_simple_neuron.x2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8468_ _4162_ _4180_ _4182_ _4183_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_103_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8399_ _3703_ ci_adder.input_memory\[1\]\[17\] _4122_ _4137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7419_ ci_adder.uut_simple_neuron.titan_id_1\[29\] ci_adder.uut_simple_neuron.titan_id_0\[29\]
+ _3437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7806__A1 _3659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8449__I3 _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5293__A1 _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8697__CLK net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5596__A2 ci_adder.uut_simple_neuron.x3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6545__A1 _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4859__A1 _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5284__A1 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4626__A4 ci_adder.uut_simple_neuron.x2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8612__I3 ci_adder.uut_simple_neuron.x3\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ _0870_ _1133_ _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7770_ ci_adder.value_i\[23\] _3629_ _3732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_106_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6721_ _1807_ _2761_ _2832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6652_ _2757_ _2763_ _2764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_85_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8525__A2 _4212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5603_ _1709_ _1715_ _1736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6583_ _2694_ _2695_ _2696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8322_ _3713_ ci_adder.uut_simple_neuron.x0\[19\] _4091_ _4094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8289__A1 _3631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5534_ _1637_ _1639_ _1672_ _1673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4562__A3 _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5465_ _1603_ _1604_ _1605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8253_ ci_adder.uut_simple_neuron.titan_id_6\[20\] _4057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5511__A2 ci_adder.uut_simple_neuron.x2\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7204_ ci_adder.uut_simple_neuron.titan_id_2\[23\] ci_adder.uut_simple_neuron.titan_id_5\[23\]
+ _3259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4416_ internal_ih.byte5\[2\] _0623_ _0632_ internal_ih.byte1\[2\] _0633_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8184_ internal_ih.spi_tx_byte_o\[4\] _3978_ _4012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5396_ _1525_ _1537_ _1538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7135_ _3201_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_70_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4347_ internal_ih.expected_byte_count\[2\] _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7066_ _3143_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8461__A1 _4165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6017_ _2103_ _2106_ _2138_ _2139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_68_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5578__A2 ci_adder.uut_simple_neuron.x3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7968_ _3765_ ci_adder.uut_simple_neuron.x2\[30\] _3840_ _3875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7811__I1 ci_adder.uut_simple_neuron.x3\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6919_ _3018_ _3020_ _3021_ _3022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7899_ internal_ih.received_byte_count\[7\] _3836_ _3837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4389__I0 internal_ih.byte4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6766__A1 _2844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8403__I _4116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5250_ _0714_ _1316_ _1356_ _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8862__CLK net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5181_ _1325_ _1327_ _1328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_3_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8940_ _0004_ net8 ci_adder.address_i\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_108_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5009__A1 ci_adder.uut_simple_neuron.x2\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8871_ _0418_ net50 ci_adder.output_memory\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8597__I2 ci_adder.uut_simple_neuron.x2\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7822_ _3770_ _3772_ _3774_ _3775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4965_ _0718_ _1058_ _1096_ _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA_fanout35_I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7753_ _3619_ _3716_ _3717_ _3718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6704_ _2814_ _2815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4841__I _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4896_ _1006_ _1012_ _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7684_ ci_adder.value_i\[9\] _3659_ _3660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6635_ _2742_ _2746_ _2747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6566_ _1756_ _2623_ _2679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5517_ _1605_ _1628_ _1560_ _1656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8305_ _3672_ _4076_ _4085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9285_ _0151_ net26 ci_adder.uut_simple_neuron.titan_id_6\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6497_ _2245_ _2364_ _2611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_100_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8521__I2 ci_adder.uut_simple_neuron.x2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8236_ _4048_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5448_ _1544_ _1546_ _1589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5496__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5379_ _1519_ _1520_ _1521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8167_ _3979_ _3995_ _3996_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7118_ ci_adder.uut_simple_neuron.titan_id_2\[8\] ci_adder.uut_simple_neuron.titan_id_5\[8\]
+ _3184_ _3185_ _3187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8098_ internal_ih.byte7\[4\] internal_ih.byte6\[4\] _3825_ _3943_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7049_ ci_adder.uut_simple_neuron.titan_id_4\[28\] ci_adder.uut_simple_neuron.titan_id_3\[28\]
+ ci_adder.uut_simple_neuron.titan_id_4\[27\] ci_adder.uut_simple_neuron.titan_id_3\[27\]
+ _3130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4471__A2 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6748__A1 _2797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8424__S _4139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4751__I _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8735__CLK net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_123_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7476__A2 _3479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6987__A1 ci_adder.uut_simple_neuron.titan_id_4\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8334__S _4091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _0813_ _0904_ _0907_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4681_ _0804_ _0841_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_83_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8587__S1 _4253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7972__I _3825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6420_ _2479_ _2481_ _2534_ _2535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_71_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4517__A3 _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6351_ ci_adder.uut_simple_neuron.x3\[20\] _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_5302_ ci_adder.uut_simple_neuron.x2\[24\] _1445_ _1446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6282_ _2353_ _2373_ _2399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7467__A2 _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9070_ _0523_ net56 ci_adder.output_val_internal\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5233_ _1371_ _1379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8021_ internal_ih.byte2\[7\] internal_ih.byte1\[7\] _3897_ _3903_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5164_ _1306_ _1302_ _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8511__S1 _4207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6978__A1 ci_adder.uut_simple_neuron.titan_id_4\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5095_ _1210_ _1211_ _1242_ _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__9190__CLK net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8019__I1 internal_ih.byte1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8923_ _0052_ net6 ci_adder.value_i\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8758__CLK net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8854_ _0401_ net19 internal_ih.current_instruction\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7805_ ci_adder.value_i\[29\] _3629_ _3761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5997_ _2119_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5402__A1 _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8785_ _0332_ net41 internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4948_ _1075_ _1100_ _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7736_ _3703_ ci_adder.uut_simple_neuron.x3\[17\] _3692_ _3704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4879_ _0992_ _0995_ _1026_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_7667_ ci_adder.uut_simple_neuron.x3\[6\] _3617_ _3646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6618_ _2669_ _2670_ _2730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7950__I0 _3723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7598_ ci_adder.uut_simple_neuron.x0\[29\] ci_adder.uut_simple_neuron.x0\[30\] _3585_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6549_ _2365_ _2475_ _2662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_104_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_9268_ _0132_ net66 ci_adder.uut_simple_neuron.titan_id_6\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9199_ _0093_ net67 ci_adder.uut_simple_neuron.titan_id_2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8219_ ci_adder.uut_simple_neuron.titan_id_6\[3\] _4040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4692__A2 ci_adder.uut_simple_neuron.x2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6969__A1 ci_adder.uut_simple_neuron.titan_id_4\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7630__A2 _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5641__A1 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7697__A2 _3629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8900__CLK net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8128__I _3811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5920_ _1995_ _2043_ _2044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5632__A1 _1735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4435__A2 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ _1935_ _1933_ _1977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_69_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5782_ _1713_ _1774_ _1908_ _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4802_ _0957_ _0942_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8570_ _4257_ _4264_ _4266_ _4267_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4733_ _0886_ _0889_ _0884_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7521_ _3519_ _3521_ _3522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_29_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7452_ _3463_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6403_ _2501_ _2503_ _2518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4664_ _0718_ _0794_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7932__I0 _3677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4595_ _0744_ _0757_ _0758_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_71_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7383_ _3403_ _3404_ _3406_ _3407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_9_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6334_ _2400_ _2437_ _2450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9122_ _0187_ net28 ci_adder.uut_simple_neuron.titan_id_0\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ _2379_ _2382_ _2383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9053_ ci_adder.input_memory\[1\]\[21\] net29 ci_adder.uut_simple_neuron.titan_id_1\[23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5216_ _1339_ _1361_ _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8004_ internal_ih.byte1\[7\] internal_ih.byte0\[7\] _3886_ _3894_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6196_ _2224_ _2315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5871__A1 ci_adder.uut_simple_neuron.x3\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5147_ _1256_ _1278_ _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5078_ ci_adder.uut_simple_neuron.x2\[18\] _1184_ _1226_ _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5623__A1 _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8906_ _0034_ net12 ci_adder.value_i\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8837_ _0384_ net15 internal_ih.byte6\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8768_ _0315_ net73 ci_adder.uut_simple_neuron.x2\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_75_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7719_ _3520_ _3682_ _3689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8699_ _0254_ net65 ci_adder.uut_simple_neuron.x3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_90_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7679__A2 _3654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8923__CLK net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_89_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5100__I _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_100_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6342__A2 _2457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4380_ internal_ih.byte4\[4\] internal_ih.byte3\[4\] _0599_ _0611_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8059__S _3919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6050_ _2122_ _2155_ _2171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_111_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5001_ _1151_ _1121_ _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_56_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Left_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6952_ ci_adder.uut_simple_neuron.titan_id_4\[12\] ci_adder.uut_simple_neuron.titan_id_3\[12\]
+ _3050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5903_ _1987_ _2007_ _2027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6883_ _2986_ _2989_ _2991_ _2992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_49_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5834_ ci_adder.uut_simple_neuron.x3\[11\] _1959_ _1960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5010__I ci_adder.uut_simple_neuron.x2\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8622_ _4166_ ci_adder.normalised_stream_write_address\[0\] _4308_ _4309_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7646__B _3599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5765_ _1834_ _1855_ _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8553_ _0697_ _4253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_8_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5696_ _1790_ _1821_ _1825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4716_ _0873_ _0874_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7504_ _3507_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8484_ ci_adder.output_memory\[7\] _4163_ _4196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4647_ _0787_ ci_adder.uut_simple_neuron.x2\[8\] _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_71_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8946__CLK net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7435_ _3449_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7366_ _3393_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6317_ _1956_ _2433_ _2434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4578_ _0714_ _0720_ _0741_ _0742_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_9105_ _0170_ net65 ci_adder.uut_simple_neuron.titan_id_0\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7297_ _3334_ _3335_ _3336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8330__I0 _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6248_ ci_adder.uut_simple_neuron.x3\[20\] _2365_ _2366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_73_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9036_ ci_adder.input_memory\[1\]\[4\] net67 ci_adder.uut_simple_neuron.titan_id_1\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5844__A1 _1947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6179_ _2100_ _2253_ _2297_ _2298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__4647__A2 ci_adder.uut_simple_neuron.x2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8633__I1 ci_adder.output_memory\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8397__I0 _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6021__A1 ci_adder.uut_simple_neuron.x3\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5835__A1 _1958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8342__S _4070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6012__A1 _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6563__A2 _2675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8969__CLK net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ _1685_ _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_26_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5481_ _1446_ _1570_ _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_53_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4501_ _0677_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4432_ _0641_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7220_ _3272_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7151_ _3214_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4363_ internal_ih.current_instruction\[1\] _0597_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6102_ _2179_ _2180_ _2183_ _2222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7082_ _3152_ _3155_ _3156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5826__A1 _1699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6033_ _2130_ _2154_ _2155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout65_I net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7984_ _3883_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6935_ ci_adder.uut_simple_neuron.titan_id_4\[9\] ci_adder.uut_simple_neuron.titan_id_3\[9\]
+ _3036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_37_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6866_ _2881_ _2917_ _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5817_ _1907_ _1909_ _1943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6797_ _1847_ _2837_ _2907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8605_ _4257_ _4292_ _4294_ _4295_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_119_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5748_ _1754_ _1846_ _1875_ _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_91_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4565__A1 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8536_ ci_adder.uut_simple_neuron.x0\[16\] ci_adder.input_memory\[1\]\[16\] ci_adder.uut_simple_neuron.x2\[16\]
+ _2098_ _4206_ _4207_ _4239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__7095__C ci_adder.uut_simple_neuron.titan_id_5\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5679_ _1692_ _1730_ _1809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_75_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8467_ ci_adder.output_val_internal\[3\] _4170_ _4183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7418_ ci_adder.uut_simple_neuron.titan_id_1\[29\] ci_adder.uut_simple_neuron.titan_id_0\[29\]
+ _3436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8398_ _4136_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9124__CLK net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7349_ ci_adder.uut_simple_neuron.titan_id_1\[17\] ci_adder.uut_simple_neuron.titan_id_0\[17\]
+ _3379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9019_ _0502_ net37 ci_adder.input_memory\[1\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__A1 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6545__A2 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4556__A1 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8298__A2 _4071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_97_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_81_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4859__A2 ci_adder.uut_simple_neuron.x2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_90_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4981_ _1109_ _1132_ _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_106_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6720_ _2190_ _2207_ _2831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6651_ _2760_ _2762_ _2763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7733__A1 _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9147__CLK net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6582_ _1750_ _2174_ _2081_ _2695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5602_ _1726_ _1728_ _1734_ _1735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__4547__A1 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5533_ _1596_ _1636_ _1672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8321_ _4093_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8289__A2 _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5464_ _1525_ _1578_ _1604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8252_ _4056_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4839__I _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5395_ _1536_ _1537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7203_ _3256_ _3257_ _3258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4415_ _0619_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8183_ ci_adder.stream_o\[28\] _3959_ _4010_ _4011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9297__CLK net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7134_ ci_adder.uut_simple_neuron.titan_id_2\[11\] ci_adder.uut_simple_neuron.titan_id_5\[11\]
+ _3200_ _3201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_1_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7065_ ci_adder.uut_simple_neuron.titan_id_4\[1\] ci_adder.uut_simple_neuron.titan_id_3\[1\]
+ _3143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6016_ _2094_ _2102_ _2138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6224__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7967_ _3874_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6918_ ci_adder.uut_simple_neuron.titan_id_4\[6\] ci_adder.uut_simple_neuron.titan_id_3\[6\]
+ ci_adder.uut_simple_neuron.titan_id_4\[5\] ci_adder.uut_simple_neuron.titan_id_3\[5\]
+ _3021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_49_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7898_ internal_ih.received_byte_count\[6\] _3834_ _3836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6849_ _2666_ _2894_ _2958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8519_ _4211_ _4222_ _4224_ _4225_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_115_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8452__A2 _4170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6463__A1 _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4529__A1 _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5180_ _1285_ _1289_ _1326_ _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_3_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8067__S _3919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__A2 ci_adder.uut_simple_neuron.x2\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwire14 _0595_ net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_8870_ _0417_ net50 ci_adder.output_memory\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8597__I3 ci_adder.uut_simple_neuron.x3\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7821_ spi_interface_cvonk.buffer\[7\] internal_ih.spi_tx_byte_o\[7\] _3773_ _3774_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_80_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4964_ _1016_ _1111_ _1087_ _1115_ _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7752_ ci_adder.value_i\[20\] _3629_ _3717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6703_ _2811_ _2813_ _2814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_fanout28_I net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4895_ _0963_ _1008_ _1048_ _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7683_ _3608_ _3659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_117_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6634_ _2364_ _2745_ _2746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6565_ _2087_ _2105_ _2678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6496_ _2593_ _2609_ _2610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5516_ _1605_ _1628_ _1655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4940__A1 _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8304_ _3667_ _4072_ _4084_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9284_ _0150_ net26 ci_adder.uut_simple_neuron.titan_id_6\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5447_ _1586_ _1587_ _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8521__I3 ci_adder.uut_simple_neuron.x3\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8235_ ci_adder.uut_simple_neuron.titan_id_6\[11\] _4048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5378_ _1400_ _1492_ _1520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8166_ internal_ih.spi_tx_byte_o\[2\] _3978_ _3996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7117_ _3186_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8097_ _3942_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7048_ _3114_ _3117_ _3128_ _3129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9312__CLK net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8999_ _0482_ net62 ci_adder.input_memory\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5184__A1 _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4931__A1 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4680_ _0830_ _0840_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6350_ _2463_ _2464_ _2465_ _2466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5301_ ci_adder.uut_simple_neuron.x2\[25\] ci_adder.uut_simple_neuron.x2\[26\] _1445_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_12_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6281_ _1699_ _2397_ _2398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5232_ _1293_ _1377_ _1378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8020_ _3902_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_114_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5163_ _1302_ _1303_ _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5094_ _1210_ _1211_ _1242_ _1243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8922_ _0051_ net10 ci_adder.value_i\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7927__A1 ci_adder.uut_simple_neuron.x2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8853_ _0400_ net19 internal_ih.current_instruction\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7804_ _3578_ _3587_ _3749_ _3760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5996_ _2073_ _2118_ _2119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8784_ _0331_ net19 internal_ih.byte0\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4947_ _1076_ _1099_ _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7735_ _3699_ _3701_ _3702_ _3703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4878_ _1032_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7666_ ci_adder.value_i\[6\] _3613_ _3644_ _3645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6617_ _2661_ _2668_ _2729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5166__A1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4913__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7950__I1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7597_ _3584_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6548_ _2468_ _2602_ _2660_ _2661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6479_ _2548_ _2550_ _2592_ _2593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9267_ _0131_ net68 ci_adder.uut_simple_neuron.titan_id_6\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9198_ _0092_ net67 ci_adder.uut_simple_neuron.titan_id_2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8218_ _4039_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8149_ _3973_ _3979_ _3980_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8702__CLK net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7918__A1 _3641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8852__CLK net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8591__A1 ci_adder.output_memory\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9208__CLK net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7909__A1 _3621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5850_ _1929_ _1932_ _1976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ _1884_ _1885_ _1908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4801_ _0934_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4732_ _0890_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7520_ _3514_ _3520_ _3521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8080__S _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4663_ _0801_ _0821_ _0823_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7451_ _3452_ _3459_ _3462_ _3463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6402_ _2513_ _2515_ _2516_ _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_114_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7932__I1 _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6896__A1 ci_adder.uut_simple_neuron.titan_id_4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4594_ _0746_ _0754_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7382_ ci_adder.uut_simple_neuron.titan_id_1\[23\] ci_adder.uut_simple_neuron.titan_id_0\[23\]
+ _3406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6333_ _1721_ _2397_ _2449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9121_ _0186_ net29 ci_adder.uut_simple_neuron.titan_id_0\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ _2380_ _2318_ _2381_ _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9052_ ci_adder.input_memory\[1\]\[20\] net36 ci_adder.uut_simple_neuron.titan_id_1\[22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5215_ _1344_ _1360_ _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8003_ _3893_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8725__CLK net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6195_ _2276_ _2313_ _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5871__A2 ci_adder.uut_simple_neuron.x3\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5146_ _1291_ _1292_ _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5077_ ci_adder.uut_simple_neuron.x2\[19\] ci_adder.uut_simple_neuron.x2\[20\] _1226_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5623__A2 _1754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8875__CLK net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8905_ _0064_ net12 ci_adder.value_i\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8836_ _0383_ net15 internal_ih.byte6\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5979_ _1960_ _2101_ _2102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_94_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8767_ _0314_ net74 ci_adder.uut_simple_neuron.x2\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_7718_ _3508_ _3687_ ci_adder.uut_simple_neuron.x0\[15\] _3688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8698_ _0253_ net83 ci_adder.uut_simple_neuron.x3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_117_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7649_ _3627_ _3628_ _3630_ _3631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_105_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9319_ _0580_ net24 ci_adder.stream_o\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5588__I _1699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7119__A2 ci_adder.uut_simple_neuron.titan_id_5\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9180__CLK net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8748__CLK net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8619__A2 _4161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _1113_ _1150_ _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__5302__A1 ci_adder.uut_simple_neuron.x2\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8898__CLK net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5605__A2 _1735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6951_ _3045_ _3047_ _3048_ _3049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_49_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5902_ _1686_ _1984_ _2026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6882_ _2900_ _2903_ _2990_ _2991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5833_ ci_adder.uut_simple_neuron.x3\[12\] ci_adder.uut_simple_neuron.x3\[13\] _1959_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_76_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8621_ _0703_ _0706_ _4308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_122_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8552_ _0698_ _4252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_118_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6581__A3 _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5764_ _1834_ _1855_ _1892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_101_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7503_ _3503_ _3506_ _3507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout10_I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5695_ _1790_ _1821_ _1823_ _1824_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4715_ ci_adder.uut_simple_neuron.x2\[9\] ci_adder.uut_simple_neuron.x2\[10\] ci_adder.uut_simple_neuron.x2\[11\]
+ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_72_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8483_ _4162_ _4192_ _4194_ _4195_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4646_ _0807_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7434_ ci_adder.uut_simple_neuron.x0\[2\] _3448_ _3449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5541__A1 ci_adder.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4577_ _0710_ _0732_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7365_ _3391_ _3392_ _3393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7530__A2 _3524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6316_ _1962_ _2432_ _2433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9104_ _0199_ net66 ci_adder.uut_simple_neuron.titan_id_0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7296_ ci_adder.uut_simple_neuron.titan_id_1\[9\] ci_adder.uut_simple_neuron.titan_id_0\[9\]
+ _3335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6247_ ci_adder.uut_simple_neuron.x3\[21\] _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_9035_ ci_adder.input_memory\[1\]\[3\] net63 ci_adder.uut_simple_neuron.titan_id_1\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_110_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6178_ _2249_ _2252_ _2297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5129_ _1119_ _1276_ _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_98_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8819_ _0366_ net16 internal_ih.byte4\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4487__I _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5835__A2 _1960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5599__A1 ci_adder.uut_simple_neuron.x3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__A2 _1958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5480_ _1611_ _1619_ _1620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4500_ internal_ih.byte3\[2\] _0670_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4431_ internal_ih.byte6\[1\] _0635_ _0632_ internal_ih.byte2\[1\] _0641_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7150_ _3212_ _3213_ _3214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4362_ _0596_ internal_ih.current_instruction\[3\] internal_ih.current_instruction\[2\]
+ _0592_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6101_ _2221_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7081_ ci_adder.uut_simple_neuron.titan_id_2\[3\] ci_adder.uut_simple_neuron.titan_id_5\[3\]
+ _3155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6032_ _2133_ _2153_ _2154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__9076__CLK net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout58_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7983_ internal_ih.byte0\[5\] internal_ih.spi_rx_byte_i\[5\] _3877_ _3883_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_124_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6934_ _3031_ _3032_ _3033_ _3034_ _3035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_119_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6865_ _2972_ _2973_ _2974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8913__CLK net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8604_ ci_adder.output_val_internal\[28\] _4161_ _4295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5816_ _1866_ _1934_ _1933_ _1942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6796_ _2240_ _2257_ _2906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5747_ _1843_ _1845_ _1875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4565__A2 ci_adder.uut_simple_neuron.x2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8535_ ci_adder.output_memory\[16\] _4212_ _4238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8000__I0 internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8466_ _4165_ _4181_ _4182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5678_ _1801_ _1807_ _1808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_75_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7417_ _3428_ _3433_ _3435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4629_ _0766_ _0769_ _0791_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8397_ _3697_ ci_adder.input_memory\[1\]\[16\] _4122_ _4136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7348_ _3378_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7279_ _3316_ _3317_ _3320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9018_ _0501_ net27 ci_adder.input_memory\[1\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_28_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8519__A1 _4211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5753__A1 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__A2 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4859__A3 ci_adder.uut_simple_neuron.x2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7321__I _3356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4492__A1 internal_ih.byte2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _1116_ _1131_ _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_106_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6650_ _1807_ _2761_ _2762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6581_ _1765_ _1796_ _1772_ _2694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5601_ _1692_ _1733_ _1734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5744__A1 _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4547__A2 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5532_ _1625_ _1665_ _1670_ _1671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_42_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8320_ _3708_ ci_adder.uut_simple_neuron.x0\[18\] _4091_ _4093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5463_ _1565_ _1577_ _1603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8251_ ci_adder.uut_simple_neuron.titan_id_6\[19\] _4056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5394_ _1528_ _1535_ _1536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7202_ _3253_ _3254_ _3257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4414_ _0631_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8182_ _3960_ _4007_ _4009_ _3815_ _4010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7133_ _3196_ _3197_ _3199_ _3200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_111_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8541__S0 _4206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7064_ _3142_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_70_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6015_ _1772_ _2136_ _2137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_68_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7966_ _3762_ ci_adder.uut_simple_neuron.x2\[29\] _3840_ _3874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6917_ _3010_ _3019_ _3020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_53_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7897_ _3826_ _3835_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6848_ _2892_ _2893_ _2957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6779_ _2887_ _2888_ _2889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8518_ ci_adder.output_val_internal\[12\] _4203_ _4225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9241__CLK net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7488__A1 ci_adder.uut_simple_neuron.x0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8449_ ci_adder.uut_simple_neuron.x0\[0\] ci_adder.input_memory\[1\]\[0\] _0710_
+ _1684_ _4166_ _4167_ _4168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_102_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6160__A1 _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8809__CLK net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8959__CLK net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7660__A1 _3608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7963__A2 _3841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5974__A1 ci_adder.uut_simple_neuron.x3\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4529__A2 _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7820_ spi_interface_cvonk.state\[2\] spi_interface_cvonk.state\[1\] spi_interface_cvonk.state\[0\]
+ _3773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_59_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9114__CLK net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5965__A1 _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4963_ _1113_ _1114_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7751_ _3539_ _3715_ _3716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6702_ ci_adder.uut_simple_neuron.x3\[26\] _2812_ _2813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7682_ _3479_ _3647_ ci_adder.uut_simple_neuron.x0\[9\] _3658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6633_ _2743_ _2744_ _2745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5717__A1 _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4894_ _0909_ _1007_ _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9264__CLK net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6564_ _2654_ _2676_ _2677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_30_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6495_ _2604_ _2608_ _2609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5515_ _1608_ _1626_ _1653_ _1654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4940__A2 ci_adder.uut_simple_neuron.x2\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8303_ ci_adder.uut_simple_neuron.x0\[10\] _4076_ _4084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9283_ _0148_ net26 ci_adder.uut_simple_neuron.titan_id_6\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5446_ _1549_ _1550_ _1585_ _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_89_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8234_ _4047_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7670__B _3470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5377_ _1477_ _1491_ _1519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7890__A1 _3826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8165_ ci_adder.stream_o\[26\] _3959_ _3994_ _3995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7116_ _3184_ _3185_ _3186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8096_ internal_ih.byte7\[3\] internal_ih.byte6\[3\] _3825_ _3942_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7047_ ci_adder.uut_simple_neuron.titan_id_4\[26\] ci_adder.uut_simple_neuron.titan_id_3\[26\]
+ _3128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4456__A1 internal_ih.byte0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_83_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7945__A2 _3841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8998_ _0481_ net62 ci_adder.input_memory\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7949_ _3865_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4931__A2 _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6133__A1 _2249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8781__CLK net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7633__A1 _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8681__I0 ci_adder.stream_o\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9137__CLK net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5300_ _0713_ _1443_ _1438_ _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6280_ _2395_ _2396_ _2397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5231_ _0994_ _1324_ _1377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8078__S _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5162_ _1304_ _1307_ _1272_ _1308_ _1234_ _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5093_ _0804_ _1241_ _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8921_ _0050_ net6 ci_adder.value_i\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8752__D _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8852_ _0399_ net19 internal_ih.current_instruction\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7927__A2 _3846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout40_I net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8783_ _0330_ net42 internal_ih.byte0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7803_ ci_adder.uut_simple_neuron.x0\[29\] _3754_ _3759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5995_ _2116_ _2117_ _2118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7734_ ci_adder.value_i\[17\] _3659_ _3702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4946_ _1078_ _1098_ _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_117_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4877_ _1029_ _1031_ _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7665_ _3613_ _3643_ _3644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6616_ _2672_ _2675_ _2727_ _2728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7596_ ci_adder.uut_simple_neuron.x0\[28\] ci_adder.uut_simple_neuron.x0\[29\] _3583_
+ _3584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6547_ _2659_ _2601_ _2660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6478_ _2542_ _2547_ _2592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_9266_ _0130_ net68 ci_adder.uut_simple_neuron.titan_id_6\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6666__A2 _2777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5429_ ci_adder.uut_simple_neuron.x2\[27\] _1530_ _1570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9197_ _0091_ net67 ci_adder.uut_simple_neuron.titan_id_2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8217_ ci_adder.uut_simple_neuron.titan_id_6\[2\] _4039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8148_ internal_ih.spi_tx_byte_o\[0\] _3979_ _3980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4429__B2 internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8079_ _3933_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_69_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5929__A1 _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7918__A2 _3841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7854__A1 internal_ih.spi_rx_byte_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6409__A2 _2496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5093__A1 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8406__I0 _3718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4840__A1 _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7909__A2 _3841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4800_ _0715_ _0932_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_14_Left_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5780_ _1694_ _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_84_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4731_ _0887_ _0889_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_83_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4662_ _0803_ _0820_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7450_ _3460_ _3461_ _3462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6401_ _2328_ _2514_ _2516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_116_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4593_ _0746_ _0754_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7705__S _3632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7381_ _3405_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9120_ _0185_ net29 ci_adder.uut_simple_neuron.titan_id_0\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6332_ _2448_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9302__CLK net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6263_ _2314_ _2317_ _2381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_86_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9051_ ci_adder.input_memory\[1\]\[19\] net36 ci_adder.uut_simple_neuron.titan_id_1\[21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_23_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5214_ _1346_ _1359_ _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8002_ internal_ih.byte1\[6\] internal_ih.byte0\[6\] _3886_ _3893_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6194_ _2278_ _2312_ _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout88_I net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5145_ _0870_ _1280_ _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5076_ _1089_ _1090_ _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8904_ _0063_ net12 ci_adder.value_i\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8835_ _0382_ net15 internal_ih.byte6\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5978_ _2097_ _2100_ _2101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8766_ _0313_ net75 ci_adder.uut_simple_neuron.x2\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7620__I1 _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4929_ _0908_ _1050_ _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8697_ _0252_ net86 ci_adder.uut_simple_neuron.x3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7717_ _3682_ _3687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7648_ ci_adder.value_i\[3\] _3629_ _3630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7579_ ci_adder.uut_simple_neuron.x0\[25\] ci_adder.uut_simple_neuron.x0\[26\] _3570_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_120_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9318_ _0579_ net24 ci_adder.stream_o\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9249_ _0114_ net72 ci_adder.uut_simple_neuron.titan_id_5\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7836__A1 internal_ih.spi_rx_byte_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4822__A1 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_100_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4889__A1 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6950_ ci_adder.uut_simple_neuron.titan_id_4\[11\] ci_adder.uut_simple_neuron.titan_id_3\[11\]
+ _3048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5066__A1 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5901_ _2023_ _2024_ _2025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4813__A1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6881_ _2886_ _2898_ _2990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6566__A1 _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5832_ ci_adder.uut_simple_neuron.x3\[10\] _1918_ _1957_ _1958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_57_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8620_ _4170_ _4304_ _4306_ _4307_ _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__8555__A2 _4254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5763_ _1867_ _1869_ _1890_ _1891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_8_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8551_ ci_adder.output_memory\[19\] _4212_ _4251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4714_ _0713_ _0854_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7502_ _3493_ _3504_ _3505_ _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5694_ _1822_ _1821_ _1824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_44_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8482_ ci_adder.output_val_internal\[6\] _4170_ _4195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4645_ _0709_ _0790_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_72_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7433_ ci_adder.uut_simple_neuron.x0\[0\] _3447_ _3448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5541__A2 _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4576_ _0740_ _0725_ _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7364_ ci_adder.uut_simple_neuron.titan_id_1\[20\] ci_adder.uut_simple_neuron.titan_id_0\[20\]
+ _3392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6315_ _2049_ _2370_ _2431_ _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9103_ _0198_ net67 ci_adder.uut_simple_neuron.titan_id_0\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7295_ _3332_ _3333_ _3334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9034_ ci_adder.input_memory\[1\]\[2\] net62 ci_adder.uut_simple_neuron.titan_id_1\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6246_ _2200_ _2301_ _2363_ _2364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__8842__CLK net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8491__A1 _4165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6177_ _2255_ _2258_ _2295_ _2296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5128_ _0811_ _1083_ _1275_ _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8992__CLK net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5059_ _1198_ _1208_ _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_43_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8818_ _0365_ net17 internal_ih.byte4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8749_ _0296_ net52 internal_ih.received_byte_count\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_23_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8537__A2 _4239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4430_ _0640_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6100_ _2218_ _2220_ _2221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4361_ internal_ih.current_instruction\[0\] _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_21_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7989__I _3825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7080_ ci_adder.uut_simple_neuron.titan_id_2\[3\] ci_adder.uut_simple_neuron.titan_id_5\[3\]
+ _3154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6031_ _2137_ _2139_ _2152_ _2153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__8086__S _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7982_ _3882_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_124_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6933_ ci_adder.uut_simple_neuron.titan_id_4\[8\] ci_adder.uut_simple_neuron.titan_id_3\[8\]
+ _3034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6864_ _1871_ _2928_ _2973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8528__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5815_ _1902_ _1938_ _1940_ _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_76_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8603_ _4260_ _4293_ _4294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_119_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6795_ _2883_ _2904_ _2905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_85_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5211__A1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5746_ _1848_ _1852_ _1873_ _1874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8534_ _4211_ _4234_ _4236_ _4237_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_115_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5677_ _1732_ _1806_ _1807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_72_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8465_ ci_adder.uut_simple_neuron.x0\[3\] ci_adder.input_memory\[1\]\[3\] _0722_
+ ci_adder.uut_simple_neuron.x3\[3\] _4166_ _4167_ _4181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_45_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8000__I1 internal_ih.byte0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4628_ _0709_ _0788_ _0790_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7416_ _3434_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8396_ _4135_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4559_ _0723_ _0725_ _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7347_ _3375_ _3377_ _3378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7278_ ci_adder.uut_simple_neuron.titan_id_1\[6\] ci_adder.uut_simple_neuron.titan_id_0\[6\]
+ _3319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8464__A1 ci_adder.output_memory\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6229_ _2345_ _2346_ _2347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9017_ _0500_ net36 ci_adder.input_memory\[1\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8067__I1 internal_ih.byte4\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9170__CLK net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5753__A2 _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6702__A1 ci_adder.uut_simple_neuron.x3\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6580_ _2691_ _2692_ _2693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5600_ _1730_ _1732_ _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5744__A2 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5531_ ci_adder.uut_simple_neuron.x2\[31\] _1668_ _1669_ _1670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_5_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8250_ _4055_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5462_ _1600_ _1601_ _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7201_ ci_adder.uut_simple_neuron.titan_id_2\[22\] ci_adder.uut_simple_neuron.titan_id_5\[22\]
+ _3256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5393_ _1482_ _1534_ _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4413_ internal_ih.byte5\[1\] _0623_ _0620_ internal_ih.byte1\[1\] _0631_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8181_ _3811_ _4008_ _4009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7132_ ci_adder.uut_simple_neuron.titan_id_2\[10\] ci_adder.uut_simple_neuron.titan_id_5\[10\]
+ _3199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7249__A2 ci_adder.uut_simple_neuron.titan_id_5\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7063_ ci_adder.uut_simple_neuron.titan_id_4\[31\] ci_adder.uut_simple_neuron.titan_id_3\[31\]
+ _3141_ _3142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8541__S1 _4207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6014_ _1778_ _2135_ _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout70_I net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9193__CLK net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4483__A2 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_6_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7965_ _3873_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6916_ _3011_ _3016_ _3019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_53_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7896_ internal_ih.received_byte_count\[6\] _3834_ _3835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_92_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6847_ _2954_ _2955_ _2956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6778_ _2601_ _2815_ _2888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5729_ _1825_ _1824_ _1857_ _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_45_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8517_ _4214_ _4223_ _4224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8448_ _0697_ _4167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8379_ ci_adder.input_memory\[1\]\[7\] _4118_ _4127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8437__A1 internal_ih.spi_rx_byte_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5423__A1 _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9066__CLK net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7723__I0 _3691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8903__CLK net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4962_ _0831_ _1052_ _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7750_ _3535_ _3700_ _3715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6701_ ci_adder.uut_simple_neuron.x3\[27\] ci_adder.uut_simple_neuron.x3\[28\] _2812_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4893_ _0831_ _1045_ _1046_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_58_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7681_ _3656_ _3657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6632_ _2418_ _2537_ _2744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7708__S _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5717__A2 _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6563_ _2672_ _2675_ _2676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4640__B _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6494_ _2249_ _2607_ _2608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5514_ _1525_ _1627_ _1653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8506__I2 ci_adder.uut_simple_neuron.x2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8302_ _4083_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9282_ _0147_ net26 ci_adder.uut_simple_neuron.titan_id_6\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5445_ _1549_ _1550_ _1585_ _1586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_70_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8233_ ci_adder.uut_simple_neuron.titan_id_6\[10\] _4047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8164_ _3960_ _3991_ _3993_ _3815_ _3994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5376_ _1475_ _1493_ _1517_ _1518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7115_ ci_adder.uut_simple_neuron.titan_id_2\[8\] ci_adder.uut_simple_neuron.titan_id_5\[8\]
+ _3185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8095_ _3941_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7046_ _3113_ _3126_ _3127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7642__A2 _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5653__A1 _1723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4815__B _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8997_ _0480_ net62 ci_adder.input_memory\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7948_ _3718_ ci_adder.uut_simple_neuron.x2\[20\] _3855_ _3865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8073__I _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7158__A1 _3216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7879_ internal_ih.received_byte_count\[1\] _3822_ _3823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5708__A2 _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6381__A2 _2496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7705__I0 _3677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8926__CLK net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7633__A2 _3617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8681__I1 ci_adder.output_memory\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5644__A1 ci_adder.uut_simple_neuron.x3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_78_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5230_ _1201_ _1206_ _1375_ _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_59_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7872__A2 _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_87_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5161_ _0718_ _1270_ _1308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5092_ _1213_ _1240_ _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5635__A1 _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8094__S _3825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8920_ _0049_ net6 ci_adder.value_i\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_69_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9231__CLK net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8851_ _0398_ net19 internal_ih.current_instruction\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5994_ _2024_ _2064_ _2117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7802_ _3758_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8782_ _0329_ net18 ci_adder.uut_simple_neuron.x2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_96_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4945_ _1088_ _1097_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7733_ _3613_ _3700_ _3701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout33_I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4876_ _1030_ _0989_ _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_62_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7664_ _3469_ _3638_ _3643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_117_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6615_ _2726_ _2671_ _2727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8949__CLK net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7595_ _3581_ _3582_ _3583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6546_ _2657_ _2539_ _2658_ _2659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6477_ _2535_ _2589_ _2590_ _2551_ _2555_ _2591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_9265_ _0129_ net68 ci_adder.uut_simple_neuron.titan_id_6\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5428_ _1348_ _1445_ _1569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9196_ _0090_ net64 ci_adder.uut_simple_neuron.titan_id_2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7863__A2 internal_ih.spi_rx_byte_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8216_ _4038_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5874__A1 ci_adder.uut_simple_neuron.x3\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5359_ _0993_ _1459_ _1501_ _1502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8147_ _3978_ _3979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8078_ internal_ih.byte6\[2\] internal_ih.byte5\[2\] _3930_ _3933_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7029_ ci_adder.uut_simple_neuron.titan_id_4\[26\] ci_adder.uut_simple_neuron.titan_id_3\[26\]
+ _3113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5626__A1 _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4429__A2 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_13_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9104__CLK net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5865__A1 _1715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7811__S _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8654__I1 ci_adder.output_memory\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__A1 _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4730_ _0865_ _0864_ _0866_ _0888_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_64_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4661_ _0822_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6400_ _2066_ _2072_ _2330_ _2514_ _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7380_ _3403_ _3404_ _3405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6331_ _2442_ _2447_ _2448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_116_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4592_ _0756_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6262_ _2265_ _2267_ _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9050_ ci_adder.input_memory\[1\]\[18\] net36 ci_adder.uut_simple_neuron.titan_id_1\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6193_ _2288_ _2290_ _2311_ _2312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5213_ _1347_ _1356_ _1358_ _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8001_ _3892_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5144_ _1249_ _1279_ _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8645__I1 ci_adder.output_memory\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5075_ _1089_ _1181_ _1124_ _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__6281__A1 _1699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8903_ _0062_ net13 ci_adder.value_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8834_ _0381_ net17 internal_ih.byte6\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5977_ ci_adder.uut_simple_neuron.x3\[14\] _2099_ _2100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_4
XFILLER_0_75_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8765_ _0312_ net37 ci_adder.uut_simple_neuron.x2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_8696_ _0251_ net88 ci_adder.uut_simple_neuron.x3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4928_ _0831_ _1052_ _1080_ _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7716_ _3686_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7647_ _3608_ _3629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6336__A2 _2408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4859_ _0899_ ci_adder.uut_simple_neuron.x2\[13\] ci_adder.uut_simple_neuron.x2\[14\]
+ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__9127__CLK net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7578_ _3565_ _3561_ _3568_ _3564_ _3569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_16_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ _2640_ _2642_ _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9317_ _0578_ net22 ci_adder.stream_o\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9248_ _0113_ net71 ci_adder.uut_simple_neuron.titan_id_5\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__A1 _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9179_ _0212_ net78 ci_adder.uut_simple_neuron.titan_id_3\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6575__A2 _2687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4586__A1 _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8572__I0 ci_adder.uut_simple_neuron.x0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8324__I0 _3718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5838__A1 _1754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5900_ _2012_ _1974_ _2011_ _2024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_72_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8794__CLK net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6015__A1 _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6880_ _2987_ _2913_ _2988_ _2989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5831_ ci_adder.uut_simple_neuron.x3\[11\] ci_adder.uut_simple_neuron.x3\[12\] _1957_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7763__A1 ci_adder.uut_simple_neuron.x0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5762_ _1872_ _1889_ _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4577__A1 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8550_ _4211_ _4246_ _4248_ _4250_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_122_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4713_ _0848_ _0857_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7501_ _3497_ _3500_ _3505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5693_ _1790_ _1822_ _1821_ _1823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8481_ _4165_ _4193_ _4194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_126_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4644_ _0788_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7432_ ci_adder.uut_simple_neuron.x0\[1\] _3447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_102_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4575_ _0709_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_7363_ ci_adder.uut_simple_neuron.titan_id_1\[19\] ci_adder.uut_simple_neuron.titan_id_0\[19\]
+ _3380_ _3388_ _3390_ _3391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__8315__I0 _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6314_ _2051_ _2199_ _2431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7294_ _3329_ _3330_ _3333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9102_ _0197_ net66 ci_adder.uut_simple_neuron.titan_id_0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6245_ _2250_ ci_adder.uut_simple_neuron.x3\[20\] _2363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5829__A1 _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9033_ ci_adder.input_memory\[1\]\[1\] net61 ci_adder.uut_simple_neuron.titan_id_1\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6176_ _2247_ _2254_ _2295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5127_ _1229_ _1231_ _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5058_ _1207_ _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7754__A1 _3632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8817_ _0364_ net23 internal_ih.byte4\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_43_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8748_ _0295_ net44 internal_ih.received_byte_count\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_23_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8679_ ci_adder.stream_o\[24\] ci_adder.output_memory\[24\] _4334_ _4339_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_23_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4740__A1 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8482__A2 _4170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6245__A1 _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8617__S0 _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_51_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4360_ internal_ih.current_instruction\[3\] _0592_ _0593_ _0594_ _0595_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_111_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6030_ _2148_ _2151_ _2152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6484__A1 _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_60_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6236__A1 _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7981_ internal_ih.byte0\[4\] internal_ih.spi_rx_byte_i\[4\] _3877_ _3882_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_124_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6932_ ci_adder.uut_simple_neuron.titan_id_4\[8\] ci_adder.uut_simple_neuron.titan_id_3\[8\]
+ ci_adder.uut_simple_neuron.titan_id_4\[7\] ci_adder.uut_simple_neuron.titan_id_3\[7\]
+ _3033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_77_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6863_ _1876_ _1886_ _2972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6539__A2 _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5814_ _1903_ _1937_ _1940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8602_ ci_adder.uut_simple_neuron.x0\[28\] ci_adder.input_memory\[1\]\[28\] _1530_
+ ci_adder.uut_simple_neuron.x3\[28\] _4252_ _4253_ _4293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_9_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6794_ _2900_ _2903_ _2904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5211__A2 ci_adder.uut_simple_neuron.x2\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5745_ _1841_ _1847_ _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8533_ ci_adder.output_val_internal\[15\] _4203_ _4237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5676_ _1803_ _1805_ _1806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4970__A1 _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8464_ ci_adder.output_memory\[3\] _4163_ _4180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4627_ _0785_ _0789_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7415_ _3432_ _3433_ _3434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_5_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8395_ _3691_ ci_adder.input_memory\[1\]\[15\] _4122_ _4135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4558_ _0724_ _0722_ _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7346_ _3376_ _3377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_12_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7277_ _3318_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4489_ _0671_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6228_ _1876_ _2293_ _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9016_ _0499_ net36 ci_adder.input_memory\[1\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6159_ _2235_ _2262_ _2277_ _2278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6227__A1 _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9315__CLK net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4961__A1 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput5 net5 spi_poci_o vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6466__A1 _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8832__CLK net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8650__S _4323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4952__A1 _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5530_ _1310_ _1340_ _1333_ _1669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5461_ _1151_ _1559_ _1601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8143__A1 internal_ih.spi_rx_byte_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4412_ _0630_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7200_ _3255_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5392_ _1529_ _1533_ _1534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_50_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8180_ ci_adder.output_val_internal\[28\] ci_adder.output_val_internal\[20\] ci_adder.output_val_internal\[12\]
+ ci_adder.output_val_internal\[4\] _3964_ _3961_ _4008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_111_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7131_ _3198_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7062_ _3137_ _3139_ _3140_ _3141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6013_ _1843_ _2104_ _2134_ _2135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_fanout63_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7964_ _3757_ _1530_ _3840_ _3873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6915_ ci_adder.uut_simple_neuron.titan_id_4\[6\] ci_adder.uut_simple_neuron.titan_id_3\[6\]
+ _3018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_53_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7895_ _3826_ _3833_ _3834_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_119_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6846_ _2953_ ci_adder.uut_simple_neuron.x3\[28\] ci_adder.uut_simple_neuron.x3\[29\]
+ _2955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8382__A1 _3654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6777_ _2811_ _2813_ _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5728_ _1827_ _1831_ _1856_ _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__4943__A1 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8516_ ci_adder.uut_simple_neuron.x0\[12\] ci_adder.input_memory\[1\]\[12\] _0899_
+ ci_adder.uut_simple_neuron.x3\[12\] _4206_ _4207_ _4223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_33_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_107_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5659_ _1789_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8447_ _0698_ _4166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_60_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8378_ _3645_ _4117_ _4126_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7329_ ci_adder.uut_simple_neuron.titan_id_1\[14\] ci_adder.uut_simple_neuron.titan_id_0\[14\]
+ _3363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_5_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5120__A1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_116_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6620__A1 ci_adder.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8460__I2 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_99_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4934__A1 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_125_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7723__I1 _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7814__S _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5662__A2 _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8444__I _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4961_ _0939_ _1112_ _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6700_ _2809_ _2810_ _2811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4892_ _1005_ _1009_ _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7680_ _3479_ ci_adder.uut_simple_neuron.x0\[9\] _3647_ _3656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_117_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6631_ _2418_ _2537_ _2743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5178__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9010__CLK net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6562_ _2141_ _2674_ _2675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_89_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8301_ _3661_ ci_adder.uut_simple_neuron.x0\[9\] _4076_ _4083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6493_ _2605_ _2606_ _2607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5513_ _1612_ _1650_ _1651_ _1652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8506__I3 ci_adder.uut_simple_neuron.x3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9281_ _0146_ net32 ci_adder.uut_simple_neuron.titan_id_6\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5444_ _0996_ _1584_ _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9160__CLK net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8232_ _4046_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8163_ _3960_ _3992_ _3993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5375_ _1437_ _1495_ _1517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7114_ _3176_ _3182_ _3183_ _3184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_10_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8094_ internal_ih.byte7\[2\] internal_ih.byte6\[2\] _3825_ _3941_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7045_ _3120_ _3122_ _3126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5102__A1 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8996_ _0479_ net52 spi_interface_cvonk.state\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7947_ _3864_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7878_ _3820_ _3821_ _0587_ _3822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6829_ _2869_ _2938_ _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8107__A1 internal_ih.spi_rx_byte_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7705__I1 ci_adder.uut_simple_neuron.x3\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4392__A2 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5341__A1 ci_adder.uut_simple_neuron.x2\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5644__A2 ci_adder.uut_simple_neuron.x3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9033__CLK net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7149__A2 ci_adder.uut_simple_neuron.titan_id_5\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5580__A1 _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5160_ _1016_ _1305_ _1260_ _1262_ _1306_ _1307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5091_ _1156_ _1239_ _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5635__A2 _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8850_ _0397_ net19 internal_ih.current_instruction\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5993_ _2074_ _2115_ _2116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7801_ _3757_ ci_adder.uut_simple_neuron.x3\[28\] _3611_ _3758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8781_ _0328_ net25 ci_adder.uut_simple_neuron.x2\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _1077_ _1096_ _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7732_ _3524_ _3695_ _3700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout26_I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4875_ _0984_ _0987_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6899__A1 ci_adder.uut_simple_neuron.titan_id_4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7663_ _3612_ _3641_ _3642_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6614_ _2656_ _2726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7594_ _3576_ _3579_ _3582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6545_ _2474_ _2538_ _2658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5571__A1 _1699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7699__I0 _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9264_ _0128_ net67 ci_adder.uut_simple_neuron.titan_id_6\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6476_ _2548_ _2550_ _2590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8215_ ci_adder.uut_simple_neuron.titan_id_6\[1\] _4038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5427_ _1566_ _1567_ _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9195_ _0089_ net64 ci_adder.uut_simple_neuron.titan_id_2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5358_ _1427_ _1458_ _1501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8146_ _3975_ _3977_ _3978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8077_ _3932_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5626__A2 _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7028_ _3112_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6823__A1 _2921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5289_ _1431_ _1432_ _1433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8979_ _0462_ net33 ci_adder.uut_simple_neuron.x0\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_65_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8328__A1 ci_adder.uut_simple_neuron.x0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6332__I _2448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7790__A2 _3629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ _0801_ _0821_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5553__A1 _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6330_ _2332_ _2443_ _2446_ _2447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_116_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4591_ _0738_ _0755_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_52_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6261_ _2376_ _2378_ _2379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_86_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _2294_ _2310_ _2311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5212_ _1310_ _1311_ _1357_ _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8000_ internal_ih.byte1\[5\] internal_ih.byte0\[5\] _3886_ _3892_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5143_ _1290_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9079__CLK net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5074_ _1186_ _1187_ _1222_ _1163_ _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_8902_ _0061_ net13 ci_adder.value_i\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_48_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8833_ _0380_ net23 internal_ih.byte6\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8916__CLK net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5976_ _2050_ _2098_ _2099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_94_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8764_ _0311_ net81 ci_adder.uut_simple_neuron.x2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5792__A1 ci_adder.uut_simple_neuron.x3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4927_ _0963_ _1079_ _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8695_ _0250_ net86 ci_adder.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_7715_ _3685_ ci_adder.uut_simple_neuron.x3\[14\] _3632_ _3686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4858_ _0899_ ci_adder.uut_simple_neuron.x2\[13\] ci_adder.uut_simple_neuron.x2\[14\]
+ _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_51_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7646_ ci_adder.uut_simple_neuron.x0\[3\] _3623_ _3599_ _3628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4789_ _0845_ _0945_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_62_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7577_ ci_adder.uut_simple_neuron.x0\[24\] ci_adder.uut_simple_neuron.x0\[25\] _3568_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9316_ _0577_ net22 ci_adder.stream_o\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6528_ _2520_ _2570_ _2641_ _2642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6459_ _2449_ _2572_ _2573_ _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9247_ _0112_ net71 ci_adder.uut_simple_neuron.titan_id_5\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9178_ _0211_ net78 ci_adder.uut_simple_neuron.titan_id_3\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__A2 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8129_ internal_ih.data_pointer\[1\] _3961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_98_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4586__A2 ci_adder.uut_simple_neuron.x2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8021__I0 internal_ih.byte2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8572__I1 ci_adder.input_memory\[1\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5838__A2 _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4510__A2 _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8939__CLK net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5830_ _1805_ _1920_ _1955_ _1956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_76_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5761_ _1874_ _1888_ _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_57_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4712_ _0870_ _0859_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8480_ _3469_ ci_adder.input_memory\[1\]\[6\] _0766_ ci_adder.uut_simple_neuron.x3\[6\]
+ _4166_ _4167_ _4193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_7500_ ci_adder.uut_simple_neuron.x0\[12\] _3504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5692_ _1762_ _1788_ _1822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7431_ _3446_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4643_ _0772_ _0802_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4574_ _0727_ _0733_ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7362_ _3383_ _3389_ _3390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6313_ _2417_ _2429_ _2430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_77_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7293_ ci_adder.uut_simple_neuron.titan_id_1\[8\] ci_adder.uut_simple_neuron.titan_id_0\[8\]
+ _3332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9101_ _0196_ net64 ci_adder.uut_simple_neuron.titan_id_0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout6 net7 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5829__A2 _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6244_ _2195_ _2303_ _2361_ _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_0_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9032_ ci_adder.input_memory\[1\]\[0\] net61 ci_adder.uut_simple_neuron.titan_id_1\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6175_ _1876_ _2293_ _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5126_ _1258_ _1273_ _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5057_ _1200_ _1201_ _1206_ _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_79_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7451__A1 _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8816_ _0363_ net21 internal_ih.byte4\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8362__I _4116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5959_ _2080_ _2081_ _2082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7754__A2 _3718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8747_ _0294_ net52 internal_ih.received_byte_count\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8678_ _4338_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9244__CLK net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7629_ _3599_ _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_35_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8562__S0 _4252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7441__I ci_adder.uut_simple_neuron.x0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6245__A2 ci_adder.uut_simple_neuron.x3\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8490__I0 _3479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7442__A1 ci_adder.uut_simple_neuron.x0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8617__S1 _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6181__A1 ci_adder.uut_simple_neuron.x3\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6484__A2 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8447__I _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8383__S _4122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7433__A1 ci_adder.uut_simple_neuron.x0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7980_ _3881_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_124_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6931_ _3023_ _3028_ _3032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6862_ _2969_ _2970_ _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5747__A1 _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5813_ _1939_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8601_ ci_adder.output_memory\[28\] _4258_ _4292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6793_ _2298_ _2902_ _2903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_45_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8532_ _4214_ _4235_ _4236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5744_ _0163_ _1871_ _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_84_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5675_ ci_adder.uut_simple_neuron.x3\[7\] _1804_ _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_5_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_20_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8463_ _4162_ _4176_ _4178_ _4179_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_103_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6172__A1 _1960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4626_ ci_adder.uut_simple_neuron.x2\[2\] ci_adder.uut_simple_neuron.x2\[3\] ci_adder.uut_simple_neuron.x2\[4\]
+ ci_adder.uut_simple_neuron.x2\[5\] _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_60_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7414_ ci_adder.uut_simple_neuron.titan_id_1\[29\] ci_adder.uut_simple_neuron.titan_id_0\[29\]
+ _3433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8394_ _4134_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7345_ ci_adder.uut_simple_neuron.titan_id_1\[17\] ci_adder.uut_simple_neuron.titan_id_0\[17\]
+ _3376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4557_ ci_adder.uut_simple_neuron.x2\[2\] _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7276_ _3316_ _3317_ _3318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4488_ internal_ih.byte2\[4\] _0670_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6227_ _1882_ _2292_ _2345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9015_ _0498_ net36 ci_adder.input_memory\[1\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7672__A1 ci_adder.value_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6158_ _2238_ _2261_ _2277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5109_ _0718_ _1221_ _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6089_ _2192_ _2194_ _2209_ _2210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_68_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7727__A2 _3659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6163__A1 _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8784__CLK net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7663__A1 _3612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4477__A1 internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5977__A1 ci_adder.uut_simple_neuron.x3\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4401__A1 internal_ih.byte4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5460_ _1084_ _1558_ _1600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4411_ internal_ih.byte5\[0\] _0623_ _0620_ internal_ih.byte1\[0\] _0630_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5391_ _0712_ _1530_ _1532_ _1533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8526__S0 _4206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7130_ _3196_ _3197_ _3198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7061_ ci_adder.uut_simple_neuron.titan_id_4\[30\] ci_adder.uut_simple_neuron.titan_id_3\[30\]
+ _3140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7654__A1 ci_adder.value_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6012_ _1845_ _1958_ _2134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
.ends

