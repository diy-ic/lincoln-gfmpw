magic
tech gf180mcuD
magscale 1 5
timestamp 1701904273
<< obsm1 >>
rect 672 1538 20328 19305
<< metal2 >>
rect 4368 20600 4424 21000
rect 4704 20600 4760 21000
rect 5712 20600 5768 21000
rect 6048 20600 6104 21000
rect 7392 20600 7448 21000
rect 8064 20600 8120 21000
rect 8400 20600 8456 21000
rect 8736 20600 8792 21000
rect 9072 20600 9128 21000
rect 9408 20600 9464 21000
rect 9744 20600 9800 21000
rect 10080 20600 10136 21000
rect 10416 20600 10472 21000
rect 10752 20600 10808 21000
rect 11088 20600 11144 21000
rect 11424 20600 11480 21000
rect 11760 20600 11816 21000
rect 12096 20600 12152 21000
rect 12768 20600 12824 21000
rect 13104 20600 13160 21000
rect 13440 20600 13496 21000
rect 13776 20600 13832 21000
rect 14448 20600 14504 21000
rect 15792 20600 15848 21000
rect 16128 20600 16184 21000
rect 17136 20600 17192 21000
rect 8400 0 8456 400
rect 9072 0 9128 400
rect 10752 0 10808 400
rect 11424 0 11480 400
rect 12768 0 12824 400
rect 13104 0 13160 400
<< obsm2 >>
rect 798 20570 4338 20600
rect 4454 20570 4674 20600
rect 4790 20570 5682 20600
rect 5798 20570 6018 20600
rect 6134 20570 7362 20600
rect 7478 20570 8034 20600
rect 8150 20570 8370 20600
rect 8486 20570 8706 20600
rect 8822 20570 9042 20600
rect 9158 20570 9378 20600
rect 9494 20570 9714 20600
rect 9830 20570 10050 20600
rect 10166 20570 10386 20600
rect 10502 20570 10722 20600
rect 10838 20570 11058 20600
rect 11174 20570 11394 20600
rect 11510 20570 11730 20600
rect 11846 20570 12066 20600
rect 12182 20570 12738 20600
rect 12854 20570 13074 20600
rect 13190 20570 13410 20600
rect 13526 20570 13746 20600
rect 13862 20570 14418 20600
rect 14534 20570 15762 20600
rect 15878 20570 16098 20600
rect 16214 20570 17106 20600
rect 17222 20570 20202 20600
rect 798 430 20202 20570
rect 798 350 8370 430
rect 8486 350 9042 430
rect 9158 350 10722 430
rect 10838 350 11394 430
rect 11510 350 12738 430
rect 12854 350 13074 430
rect 13190 350 20202 430
<< metal3 >>
rect 0 18144 400 18200
rect 20600 15792 21000 15848
rect 0 15456 400 15512
rect 20600 15456 21000 15512
rect 0 15120 400 15176
rect 0 14448 400 14504
rect 20600 14448 21000 14504
rect 0 14112 400 14168
rect 20600 14112 21000 14168
rect 0 12768 400 12824
rect 20600 12768 21000 12824
rect 0 12432 400 12488
rect 20600 12432 21000 12488
rect 0 12096 400 12152
rect 0 11760 400 11816
rect 20600 11760 21000 11816
rect 0 11424 400 11480
rect 20600 11424 21000 11480
rect 0 11088 400 11144
rect 20600 11088 21000 11144
rect 0 10752 400 10808
rect 20600 10752 21000 10808
rect 0 10416 400 10472
rect 20600 10416 21000 10472
rect 0 10080 400 10136
rect 20600 10080 21000 10136
rect 0 9744 400 9800
rect 20600 9744 21000 9800
rect 0 9408 400 9464
rect 20600 9408 21000 9464
rect 0 9072 400 9128
rect 0 8736 400 8792
rect 0 8400 400 8456
rect 20600 8400 21000 8456
rect 0 8064 400 8120
rect 20600 8064 21000 8120
rect 0 7728 400 7784
rect 20600 7728 21000 7784
rect 20600 7392 21000 7448
rect 20600 7056 21000 7112
rect 20600 6720 21000 6776
rect 20600 6384 21000 6440
<< obsm3 >>
rect 400 18230 20600 19306
rect 430 18114 20600 18230
rect 400 15878 20600 18114
rect 400 15762 20570 15878
rect 400 15542 20600 15762
rect 430 15426 20570 15542
rect 400 15206 20600 15426
rect 430 15090 20600 15206
rect 400 14534 20600 15090
rect 430 14418 20570 14534
rect 400 14198 20600 14418
rect 430 14082 20570 14198
rect 400 12854 20600 14082
rect 430 12738 20570 12854
rect 400 12518 20600 12738
rect 430 12402 20570 12518
rect 400 12182 20600 12402
rect 430 12066 20600 12182
rect 400 11846 20600 12066
rect 430 11730 20570 11846
rect 400 11510 20600 11730
rect 430 11394 20570 11510
rect 400 11174 20600 11394
rect 430 11058 20570 11174
rect 400 10838 20600 11058
rect 430 10722 20570 10838
rect 400 10502 20600 10722
rect 430 10386 20570 10502
rect 400 10166 20600 10386
rect 430 10050 20570 10166
rect 400 9830 20600 10050
rect 430 9714 20570 9830
rect 400 9494 20600 9714
rect 430 9378 20570 9494
rect 400 9158 20600 9378
rect 430 9042 20600 9158
rect 400 8822 20600 9042
rect 430 8706 20600 8822
rect 400 8486 20600 8706
rect 430 8370 20570 8486
rect 400 8150 20600 8370
rect 430 8034 20570 8150
rect 400 7814 20600 8034
rect 430 7698 20570 7814
rect 400 7478 20600 7698
rect 400 7362 20570 7478
rect 400 7142 20600 7362
rect 400 7026 20570 7142
rect 400 6806 20600 7026
rect 400 6690 20570 6806
rect 400 6470 20600 6690
rect 400 6354 20570 6470
rect 400 1554 20600 6354
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< labels >>
rlabel metal3 s 0 18144 400 18200 6 clock
port 1 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 logisim_clock_tree_0_out
port 2 nsew signal output
rlabel metal3 s 20600 8400 21000 8456 6 ram_addr_o[0]
port 3 nsew signal output
rlabel metal3 s 20600 8064 21000 8120 6 ram_addr_o[1]
port 4 nsew signal output
rlabel metal3 s 20600 7728 21000 7784 6 ram_addr_o[2]
port 5 nsew signal output
rlabel metal2 s 13104 0 13160 400 6 ram_addr_o[3]
port 6 nsew signal output
rlabel metal3 s 20600 7392 21000 7448 6 ram_addr_o[4]
port 7 nsew signal output
rlabel metal3 s 20600 7056 21000 7112 6 ram_data_i[0]
port 8 nsew signal input
rlabel metal3 s 0 8736 400 8792 6 ram_data_i[10]
port 9 nsew signal input
rlabel metal3 s 0 9072 400 9128 6 ram_data_i[11]
port 10 nsew signal input
rlabel metal3 s 0 11088 400 11144 6 ram_data_i[12]
port 11 nsew signal input
rlabel metal3 s 0 8400 400 8456 6 ram_data_i[13]
port 12 nsew signal input
rlabel metal3 s 0 12096 400 12152 6 ram_data_i[14]
port 13 nsew signal input
rlabel metal3 s 0 11760 400 11816 6 ram_data_i[15]
port 14 nsew signal input
rlabel metal3 s 0 14448 400 14504 6 ram_data_i[16]
port 15 nsew signal input
rlabel metal3 s 0 15456 400 15512 6 ram_data_i[17]
port 16 nsew signal input
rlabel metal2 s 4704 20600 4760 21000 6 ram_data_i[18]
port 17 nsew signal input
rlabel metal2 s 5712 20600 5768 21000 6 ram_data_i[19]
port 18 nsew signal input
rlabel metal3 s 20600 6384 21000 6440 6 ram_data_i[1]
port 19 nsew signal input
rlabel metal2 s 8736 20600 8792 21000 6 ram_data_i[20]
port 20 nsew signal input
rlabel metal2 s 8400 20600 8456 21000 6 ram_data_i[21]
port 21 nsew signal input
rlabel metal2 s 9072 20600 9128 21000 6 ram_data_i[22]
port 22 nsew signal input
rlabel metal2 s 9408 20600 9464 21000 6 ram_data_i[23]
port 23 nsew signal input
rlabel metal2 s 11088 20600 11144 21000 6 ram_data_i[24]
port 24 nsew signal input
rlabel metal2 s 11760 20600 11816 21000 6 ram_data_i[25]
port 25 nsew signal input
rlabel metal2 s 13440 20600 13496 21000 6 ram_data_i[26]
port 26 nsew signal input
rlabel metal2 s 13776 20600 13832 21000 6 ram_data_i[27]
port 27 nsew signal input
rlabel metal2 s 15792 20600 15848 21000 6 ram_data_i[28]
port 28 nsew signal input
rlabel metal3 s 20600 15792 21000 15848 6 ram_data_i[29]
port 29 nsew signal input
rlabel metal3 s 20600 10080 21000 10136 6 ram_data_i[2]
port 30 nsew signal input
rlabel metal3 s 20600 15456 21000 15512 6 ram_data_i[30]
port 31 nsew signal input
rlabel metal3 s 20600 14112 21000 14168 6 ram_data_i[31]
port 32 nsew signal input
rlabel metal3 s 20600 9408 21000 9464 6 ram_data_i[3]
port 33 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 ram_data_i[4]
port 34 nsew signal input
rlabel metal3 s 20600 10752 21000 10808 6 ram_data_i[5]
port 35 nsew signal input
rlabel metal2 s 10752 20600 10808 21000 6 ram_data_i[6]
port 36 nsew signal input
rlabel metal3 s 20600 11424 21000 11480 6 ram_data_i[7]
port 37 nsew signal input
rlabel metal3 s 0 10416 400 10472 6 ram_data_i[8]
port 38 nsew signal input
rlabel metal3 s 0 10080 400 10136 6 ram_data_i[9]
port 39 nsew signal input
rlabel metal3 s 20600 11088 21000 11144 6 ram_data_o[0]
port 40 nsew signal output
rlabel metal3 s 0 7728 400 7784 6 ram_data_o[10]
port 41 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 ram_data_o[11]
port 42 nsew signal output
rlabel metal3 s 0 10752 400 10808 6 ram_data_o[12]
port 43 nsew signal output
rlabel metal3 s 0 9408 400 9464 6 ram_data_o[13]
port 44 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 ram_data_o[14]
port 45 nsew signal output
rlabel metal3 s 0 12432 400 12488 6 ram_data_o[15]
port 46 nsew signal output
rlabel metal3 s 0 14112 400 14168 6 ram_data_o[16]
port 47 nsew signal output
rlabel metal3 s 0 15120 400 15176 6 ram_data_o[17]
port 48 nsew signal output
rlabel metal2 s 4368 20600 4424 21000 6 ram_data_o[18]
port 49 nsew signal output
rlabel metal2 s 6048 20600 6104 21000 6 ram_data_o[19]
port 50 nsew signal output
rlabel metal3 s 20600 9744 21000 9800 6 ram_data_o[1]
port 51 nsew signal output
rlabel metal2 s 9744 20600 9800 21000 6 ram_data_o[20]
port 52 nsew signal output
rlabel metal2 s 7392 20600 7448 21000 6 ram_data_o[21]
port 53 nsew signal output
rlabel metal2 s 8064 20600 8120 21000 6 ram_data_o[22]
port 54 nsew signal output
rlabel metal2 s 10416 20600 10472 21000 6 ram_data_o[23]
port 55 nsew signal output
rlabel metal2 s 11424 20600 11480 21000 6 ram_data_o[24]
port 56 nsew signal output
rlabel metal2 s 12768 20600 12824 21000 6 ram_data_o[25]
port 57 nsew signal output
rlabel metal2 s 14448 20600 14504 21000 6 ram_data_o[26]
port 58 nsew signal output
rlabel metal2 s 13104 20600 13160 21000 6 ram_data_o[27]
port 59 nsew signal output
rlabel metal2 s 17136 20600 17192 21000 6 ram_data_o[28]
port 60 nsew signal output
rlabel metal2 s 16128 20600 16184 21000 6 ram_data_o[29]
port 61 nsew signal output
rlabel metal3 s 20600 12768 21000 12824 6 ram_data_o[2]
port 62 nsew signal output
rlabel metal3 s 20600 14448 21000 14504 6 ram_data_o[30]
port 63 nsew signal output
rlabel metal3 s 20600 6720 21000 6776 6 ram_data_o[31]
port 64 nsew signal output
rlabel metal3 s 20600 12432 21000 12488 6 ram_data_o[3]
port 65 nsew signal output
rlabel metal3 s 20600 11760 21000 11816 6 ram_data_o[4]
port 66 nsew signal output
rlabel metal3 s 20600 10416 21000 10472 6 ram_data_o[5]
port 67 nsew signal output
rlabel metal2 s 10080 20600 10136 21000 6 ram_data_o[6]
port 68 nsew signal output
rlabel metal2 s 12096 20600 12152 21000 6 ram_data_o[7]
port 69 nsew signal output
rlabel metal3 s 0 11424 400 11480 6 ram_data_o[8]
port 70 nsew signal output
rlabel metal3 s 0 9744 400 9800 6 ram_data_o[9]
port 71 nsew signal output
rlabel metal2 s 10752 0 10808 400 6 ram_rw_en_o
port 72 nsew signal output
rlabel metal2 s 11424 0 11480 400 6 reset_i
port 73 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 stop_lamp_o
port 74 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 75 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 75 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 76 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1568720
string GDS_FILE /home/kris/repos/diy-ic/lincoln-gfmpw/openlane/manchester-baby/runs/23_12_06_23_08/results/signoff/manchester_baby.magic.gds
string GDS_START 366846
<< end >>

