/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : main                                                         **
 **                                                                          **
 *****************************************************************************/

module main( A,
             ADC,
             AND,
             ASL,
             BCC,
             BCS,
             BEQ,
             BMI,
             BNE,
             BPL,
             BRK,
             BVC,
             BVS,
             CLC,
             CLD,
             CLI,
             CLV,
             CMP,
             CPX,
             CPY,
             DEC,
             DES,
             DEY,
             EOR,
             INC,
             INX,
             INY,
             JMP,
             JSR,
             LDA,
             LDX,
             LDX_Y,
             LDY,
             LSR,
             ORA,
             PHA,
             PHP,
             PLA,
             PLP,
             ROL,
             ROR,
             RTI,
             RTS,
             SBC,
             SEC,
             SED,
             SEI,
             STA,
             STX,
             STY,
             TAX,
             TAY,
             TKA,
             TKS,
             TSX,
             TYA,
             Xind,
             abs,
             absX,
             absY,
             hash,
             ind,
             indY,
             instruction_bus,
             rel,
             zpg,
             zpgX );

   /*******************************************************************************
   ** The inputs are defined here                                                **
   *******************************************************************************/
   input [7:0] instruction_bus;

   /*******************************************************************************
   ** The outputs are defined here                                               **
   *******************************************************************************/
   output A;
   output ADC;
   output AND;
   output ASL;
   output BCC;
   output BCS;
   output BEQ;
   output BMI;
   output BNE;
   output BPL;
   output BRK;
   output BVC;
   output BVS;
   output CLC;
   output CLD;
   output CLI;
   output CLV;
   output CMP;
   output CPX;
   output CPY;
   output DEC;
   output DES;
   output DEY;
   output EOR;
   output INC;
   output INX;
   output INY;
   output JMP;
   output JSR;
   output LDA;
   output LDX;
   output LDX_Y;
   output LDY;
   output LSR;
   output ORA;
   output PHA;
   output PHP;
   output PLA;
   output PLP;
   output ROL;
   output ROR;
   output RTI;
   output RTS;
   output SBC;
   output SEC;
   output SED;
   output SEI;
   output STA;
   output STX;
   output STY;
   output TAX;
   output TAY;
   output TKA;
   output TKS;
   output TSX;
   output TYA;
   output Xind;
   output abs;
   output absX;
   output absY;
   output hash;
   output ind;
   output indY;
   output rel;
   output zpg;
   output zpgX;

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire [7:0] s_logisimBus100;
   wire       s_logisimNet0;
   wire       s_logisimNet1;
   wire       s_logisimNet10;
   wire       s_logisimNet101;
   wire       s_logisimNet102;
   wire       s_logisimNet103;
   wire       s_logisimNet104;
   wire       s_logisimNet105;
   wire       s_logisimNet106;
   wire       s_logisimNet107;
   wire       s_logisimNet108;
   wire       s_logisimNet109;
   wire       s_logisimNet11;
   wire       s_logisimNet110;
   wire       s_logisimNet111;
   wire       s_logisimNet112;
   wire       s_logisimNet113;
   wire       s_logisimNet114;
   wire       s_logisimNet115;
   wire       s_logisimNet116;
   wire       s_logisimNet117;
   wire       s_logisimNet118;
   wire       s_logisimNet119;
   wire       s_logisimNet12;
   wire       s_logisimNet120;
   wire       s_logisimNet121;
   wire       s_logisimNet122;
   wire       s_logisimNet123;
   wire       s_logisimNet124;
   wire       s_logisimNet125;
   wire       s_logisimNet126;
   wire       s_logisimNet127;
   wire       s_logisimNet128;
   wire       s_logisimNet129;
   wire       s_logisimNet13;
   wire       s_logisimNet130;
   wire       s_logisimNet131;
   wire       s_logisimNet132;
   wire       s_logisimNet133;
   wire       s_logisimNet134;
   wire       s_logisimNet135;
   wire       s_logisimNet137;
   wire       s_logisimNet138;
   wire       s_logisimNet139;
   wire       s_logisimNet14;
   wire       s_logisimNet140;
   wire       s_logisimNet141;
   wire       s_logisimNet142;
   wire       s_logisimNet143;
   wire       s_logisimNet144;
   wire       s_logisimNet145;
   wire       s_logisimNet146;
   wire       s_logisimNet147;
   wire       s_logisimNet148;
   wire       s_logisimNet149;
   wire       s_logisimNet15;
   wire       s_logisimNet150;
   wire       s_logisimNet151;
   wire       s_logisimNet152;
   wire       s_logisimNet153;
   wire       s_logisimNet154;
   wire       s_logisimNet155;
   wire       s_logisimNet156;
   wire       s_logisimNet157;
   wire       s_logisimNet158;
   wire       s_logisimNet159;
   wire       s_logisimNet16;
   wire       s_logisimNet160;
   wire       s_logisimNet161;
   wire       s_logisimNet162;
   wire       s_logisimNet163;
   wire       s_logisimNet164;
   wire       s_logisimNet165;
   wire       s_logisimNet166;
   wire       s_logisimNet167;
   wire       s_logisimNet168;
   wire       s_logisimNet169;
   wire       s_logisimNet17;
   wire       s_logisimNet170;
   wire       s_logisimNet171;
   wire       s_logisimNet172;
   wire       s_logisimNet173;
   wire       s_logisimNet174;
   wire       s_logisimNet175;
   wire       s_logisimNet176;
   wire       s_logisimNet177;
   wire       s_logisimNet178;
   wire       s_logisimNet179;
   wire       s_logisimNet18;
   wire       s_logisimNet180;
   wire       s_logisimNet181;
   wire       s_logisimNet182;
   wire       s_logisimNet183;
   wire       s_logisimNet184;
   wire       s_logisimNet185;
   wire       s_logisimNet186;
   wire       s_logisimNet187;
   wire       s_logisimNet188;
   wire       s_logisimNet189;
   wire       s_logisimNet19;
   wire       s_logisimNet190;
   wire       s_logisimNet191;
   wire       s_logisimNet192;
   wire       s_logisimNet193;
   wire       s_logisimNet194;
   wire       s_logisimNet195;
   wire       s_logisimNet196;
   wire       s_logisimNet197;
   wire       s_logisimNet198;
   wire       s_logisimNet199;
   wire       s_logisimNet2;
   wire       s_logisimNet20;
   wire       s_logisimNet200;
   wire       s_logisimNet201;
   wire       s_logisimNet202;
   wire       s_logisimNet203;
   wire       s_logisimNet204;
   wire       s_logisimNet205;
   wire       s_logisimNet206;
   wire       s_logisimNet207;
   wire       s_logisimNet208;
   wire       s_logisimNet209;
   wire       s_logisimNet21;
   wire       s_logisimNet210;
   wire       s_logisimNet211;
   wire       s_logisimNet212;
   wire       s_logisimNet213;
   wire       s_logisimNet214;
   wire       s_logisimNet215;
   wire       s_logisimNet216;
   wire       s_logisimNet217;
   wire       s_logisimNet218;
   wire       s_logisimNet219;
   wire       s_logisimNet22;
   wire       s_logisimNet220;
   wire       s_logisimNet221;
   wire       s_logisimNet222;
   wire       s_logisimNet223;
   wire       s_logisimNet224;
   wire       s_logisimNet225;
   wire       s_logisimNet226;
   wire       s_logisimNet227;
   wire       s_logisimNet228;
   wire       s_logisimNet229;
   wire       s_logisimNet23;
   wire       s_logisimNet230;
   wire       s_logisimNet231;
   wire       s_logisimNet232;
   wire       s_logisimNet233;
   wire       s_logisimNet234;
   wire       s_logisimNet235;
   wire       s_logisimNet236;
   wire       s_logisimNet237;
   wire       s_logisimNet238;
   wire       s_logisimNet239;
   wire       s_logisimNet24;
   wire       s_logisimNet240;
   wire       s_logisimNet241;
   wire       s_logisimNet242;
   wire       s_logisimNet243;
   wire       s_logisimNet244;
   wire       s_logisimNet245;
   wire       s_logisimNet246;
   wire       s_logisimNet247;
   wire       s_logisimNet248;
   wire       s_logisimNet249;
   wire       s_logisimNet25;
   wire       s_logisimNet250;
   wire       s_logisimNet251;
   wire       s_logisimNet252;
   wire       s_logisimNet253;
   wire       s_logisimNet254;
   wire       s_logisimNet255;
   wire       s_logisimNet256;
   wire       s_logisimNet257;
   wire       s_logisimNet258;
   wire       s_logisimNet259;
   wire       s_logisimNet26;
   wire       s_logisimNet260;
   wire       s_logisimNet261;
   wire       s_logisimNet262;
   wire       s_logisimNet263;
   wire       s_logisimNet264;
   wire       s_logisimNet265;
   wire       s_logisimNet266;
   wire       s_logisimNet267;
   wire       s_logisimNet268;
   wire       s_logisimNet269;
   wire       s_logisimNet27;
   wire       s_logisimNet270;
   wire       s_logisimNet271;
   wire       s_logisimNet272;
   wire       s_logisimNet273;
   wire       s_logisimNet274;
   wire       s_logisimNet275;
   wire       s_logisimNet276;
   wire       s_logisimNet277;
   wire       s_logisimNet278;
   wire       s_logisimNet279;
   wire       s_logisimNet28;
   wire       s_logisimNet280;
   wire       s_logisimNet281;
   wire       s_logisimNet282;
   wire       s_logisimNet283;
   wire       s_logisimNet284;
   wire       s_logisimNet285;
   wire       s_logisimNet286;
   wire       s_logisimNet287;
   wire       s_logisimNet288;
   wire       s_logisimNet289;
   wire       s_logisimNet29;
   wire       s_logisimNet290;
   wire       s_logisimNet291;
   wire       s_logisimNet292;
   wire       s_logisimNet293;
   wire       s_logisimNet294;
   wire       s_logisimNet295;
   wire       s_logisimNet296;
   wire       s_logisimNet297;
   wire       s_logisimNet298;
   wire       s_logisimNet299;
   wire       s_logisimNet3;
   wire       s_logisimNet30;
   wire       s_logisimNet300;
   wire       s_logisimNet301;
   wire       s_logisimNet302;
   wire       s_logisimNet303;
   wire       s_logisimNet304;
   wire       s_logisimNet305;
   wire       s_logisimNet306;
   wire       s_logisimNet307;
   wire       s_logisimNet308;
   wire       s_logisimNet309;
   wire       s_logisimNet31;
   wire       s_logisimNet310;
   wire       s_logisimNet311;
   wire       s_logisimNet312;
   wire       s_logisimNet313;
   wire       s_logisimNet314;
   wire       s_logisimNet315;
   wire       s_logisimNet316;
   wire       s_logisimNet317;
   wire       s_logisimNet318;
   wire       s_logisimNet319;
   wire       s_logisimNet32;
   wire       s_logisimNet320;
   wire       s_logisimNet321;
   wire       s_logisimNet322;
   wire       s_logisimNet323;
   wire       s_logisimNet324;
   wire       s_logisimNet325;
   wire       s_logisimNet326;
   wire       s_logisimNet327;
   wire       s_logisimNet328;
   wire       s_logisimNet329;
   wire       s_logisimNet33;
   wire       s_logisimNet330;
   wire       s_logisimNet331;
   wire       s_logisimNet332;
   wire       s_logisimNet333;
   wire       s_logisimNet334;
   wire       s_logisimNet335;
   wire       s_logisimNet336;
   wire       s_logisimNet337;
   wire       s_logisimNet338;
   wire       s_logisimNet339;
   wire       s_logisimNet34;
   wire       s_logisimNet340;
   wire       s_logisimNet341;
   wire       s_logisimNet342;
   wire       s_logisimNet343;
   wire       s_logisimNet344;
   wire       s_logisimNet345;
   wire       s_logisimNet346;
   wire       s_logisimNet347;
   wire       s_logisimNet348;
   wire       s_logisimNet349;
   wire       s_logisimNet35;
   wire       s_logisimNet350;
   wire       s_logisimNet351;
   wire       s_logisimNet352;
   wire       s_logisimNet353;
   wire       s_logisimNet354;
   wire       s_logisimNet355;
   wire       s_logisimNet356;
   wire       s_logisimNet357;
   wire       s_logisimNet358;
   wire       s_logisimNet359;
   wire       s_logisimNet36;
   wire       s_logisimNet360;
   wire       s_logisimNet361;
   wire       s_logisimNet362;
   wire       s_logisimNet363;
   wire       s_logisimNet364;
   wire       s_logisimNet365;
   wire       s_logisimNet366;
   wire       s_logisimNet367;
   wire       s_logisimNet368;
   wire       s_logisimNet369;
   wire       s_logisimNet37;
   wire       s_logisimNet370;
   wire       s_logisimNet371;
   wire       s_logisimNet372;
   wire       s_logisimNet373;
   wire       s_logisimNet374;
   wire       s_logisimNet375;
   wire       s_logisimNet376;
   wire       s_logisimNet377;
   wire       s_logisimNet378;
   wire       s_logisimNet379;
   wire       s_logisimNet38;
   wire       s_logisimNet380;
   wire       s_logisimNet381;
   wire       s_logisimNet382;
   wire       s_logisimNet39;
   wire       s_logisimNet4;
   wire       s_logisimNet40;
   wire       s_logisimNet41;
   wire       s_logisimNet42;
   wire       s_logisimNet43;
   wire       s_logisimNet44;
   wire       s_logisimNet45;
   wire       s_logisimNet46;
   wire       s_logisimNet47;
   wire       s_logisimNet48;
   wire       s_logisimNet49;
   wire       s_logisimNet5;
   wire       s_logisimNet50;
   wire       s_logisimNet51;
   wire       s_logisimNet52;
   wire       s_logisimNet53;
   wire       s_logisimNet54;
   wire       s_logisimNet55;
   wire       s_logisimNet56;
   wire       s_logisimNet57;
   wire       s_logisimNet58;
   wire       s_logisimNet59;
   wire       s_logisimNet6;
   wire       s_logisimNet60;
   wire       s_logisimNet61;
   wire       s_logisimNet62;
   wire       s_logisimNet63;
   wire       s_logisimNet64;
   wire       s_logisimNet65;
   wire       s_logisimNet66;
   wire       s_logisimNet67;
   wire       s_logisimNet68;
   wire       s_logisimNet69;
   wire       s_logisimNet7;
   wire       s_logisimNet70;
   wire       s_logisimNet71;
   wire       s_logisimNet72;
   wire       s_logisimNet73;
   wire       s_logisimNet74;
   wire       s_logisimNet75;
   wire       s_logisimNet76;
   wire       s_logisimNet77;
   wire       s_logisimNet78;
   wire       s_logisimNet79;
   wire       s_logisimNet8;
   wire       s_logisimNet80;
   wire       s_logisimNet81;
   wire       s_logisimNet82;
   wire       s_logisimNet83;
   wire       s_logisimNet84;
   wire       s_logisimNet85;
   wire       s_logisimNet86;
   wire       s_logisimNet87;
   wire       s_logisimNet88;
   wire       s_logisimNet89;
   wire       s_logisimNet9;
   wire       s_logisimNet90;
   wire       s_logisimNet91;
   wire       s_logisimNet92;
   wire       s_logisimNet93;
   wire       s_logisimNet95;
   wire       s_logisimNet96;
   wire       s_logisimNet97;
   wire       s_logisimNet98;
   wire       s_logisimNet99;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** Here all input connections are defined                                     **
   *******************************************************************************/
   assign s_logisimBus100[7:0] = instruction_bus;

   /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
   assign A     = s_logisimNet155;
   assign ADC   = s_logisimNet28;
   assign AND   = s_logisimNet325;
   assign ASL   = s_logisimNet110;
   assign BCC   = s_logisimNet152;
   assign BCS   = s_logisimNet188;
   assign BEQ   = s_logisimNet137;
   assign BMI   = s_logisimNet82;
   assign BNE   = s_logisimNet223;
   assign BPL   = s_logisimNet51;
   assign BRK   = s_logisimNet311;
   assign BVC   = s_logisimNet222;
   assign BVS   = s_logisimNet35;
   assign CLC   = s_logisimNet302;
   assign CLD   = s_logisimNet368;
   assign CLI   = s_logisimNet367;
   assign CLV   = s_logisimNet303;
   assign CMP   = s_logisimNet330;
   assign CPX   = s_logisimNet151;
   assign CPY   = s_logisimNet294;
   assign DEC   = s_logisimNet78;
   assign DES   = s_logisimNet349;
   assign DEY   = s_logisimNet298;
   assign EOR   = s_logisimNet357;
   assign INC   = s_logisimNet180;
   assign INX   = s_logisimNet262;
   assign INY   = s_logisimNet379;
   assign JMP   = s_logisimNet382;
   assign JSR   = s_logisimNet160;
   assign LDA   = s_logisimNet189;
   assign LDX   = s_logisimNet125;
   assign LDX_Y = s_logisimNet161;
   assign LDY   = s_logisimNet124;
   assign LSR   = s_logisimNet76;
   assign ORA   = s_logisimNet121;
   assign PHA   = s_logisimNet66;
   assign PHP   = s_logisimNet359;
   assign PLA   = s_logisimNet219;
   assign PLP   = s_logisimNet372;
   assign ROL   = s_logisimNet191;
   assign ROR   = s_logisimNet11;
   assign RTI   = s_logisimNet370;
   assign RTS   = s_logisimNet380;
   assign SBC   = s_logisimNet63;
   assign SEC   = s_logisimNet340;
   assign SED   = s_logisimNet115;
   assign SEI   = s_logisimNet374;
   assign STA   = s_logisimNet327;
   assign STX   = s_logisimNet337;
   assign STY   = s_logisimNet30;
   assign TAX   = s_logisimNet258;
   assign TAY   = s_logisimNet352;
   assign TKA   = s_logisimNet62;
   assign TKS   = s_logisimNet365;
   assign TSX   = s_logisimNet112;
   assign TYA   = s_logisimNet127;
   assign Xind  = s_logisimNet378;
   assign abs   = s_logisimNet354;
   assign absX  = s_logisimNet200;
   assign absY  = s_logisimNet285;
   assign hash  = s_logisimNet371;
   assign ind   = s_logisimNet176;
   assign indY  = s_logisimNet324;
   assign rel   = s_logisimNet267;
   assign zpg   = s_logisimNet308;
   assign zpgX  = s_logisimNet363;

   /*******************************************************************************
   ** Here all normal components are defined                                     **
   *******************************************************************************/
   AND_GATE #(.BubblesMask(2'b00))
      GATES_1 (.input1(s_logisimNet85),
               .input2(s_logisimNet64),
               .result(s_logisimNet192));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_2 (.input1(s_logisimNet26),
               .input2(s_logisimNet64),
               .result(s_logisimNet271));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_3 (.input1(s_logisimNet17),
               .input2(s_logisimNet0),
               .result(s_logisimNet93));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_4 (.input1(s_logisimNet103),
               .input2(s_logisimNet305),
               .result(s_logisimNet63));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_5 (.input1(s_logisimNet27),
               .input2(s_logisimNet102),
               .result(s_logisimNet105));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_6 (.input1(s_logisimNet255),
               .input2(s_logisimNet226),
               .result(s_logisimNet323));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_7 (.input1(s_logisimNet56),
               .input2(s_logisimNet89),
               .result(s_logisimNet226));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_8 (.input1(s_logisimNet149),
               .input2(s_logisimNet7),
               .result(s_logisimNet112));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_9 (.input1(s_logisimNet85),
               .input2(s_logisimNet7),
               .result(s_logisimNet25));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_10 (.input1(s_logisimNet313),
                .input2(s_logisimNet42),
                .result(s_logisimNet234));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_11 (.input1(s_logisimNet53),
                .input2(s_logisimNet32),
                .result(s_logisimNet68));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_12 (.input1(s_logisimNet27),
                .input2(s_logisimNet29),
                .result(s_logisimNet361));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_13 (.input1(s_logisimNet111),
                .input2(s_logisimNet229),
                .result(s_logisimNet76));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_14 (.input1(s_logisimNet33),
                .input2(s_logisimNet213),
                .result(s_logisimNet206));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_15 (.input1(s_logisimNet106),
                .input2(s_logisimNet81),
                .result(s_logisimNet55));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_16 (.input1(s_logisimNet35),
                .input2(s_logisimNet235),
                .result(s_logisimNet101));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_17 (.input1(s_logisimNet74),
                .input2(s_logisimNet1),
                .result(s_logisimNet207));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_18 (.input1(s_logisimNet218),
                .input2(s_logisimNet316),
                .result(s_logisimNet377));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_19 (.input1(s_logisimNet85),
                .input2(s_logisimNet0),
                .result(s_logisimNet80));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_20 (.input1(s_logisimNet113),
                .input2(s_logisimNet287),
                .result(s_logisimNet228));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_21 (.input1(s_logisimNet75),
                .input2(s_logisimNet0),
                .result(s_logisimNet10));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_22 (.input1(s_logisimNet97),
                .input2(s_logisimNet118),
                .result(s_logisimNet244));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_23 (.input1(s_logisimNet290),
                .input2(s_logisimNet299),
                .result(s_logisimNet326));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_24 (.input1(s_logisimNet82),
                .input2(s_logisimNet51),
                .result(s_logisimNet108));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_25 (.input1(s_logisimNet93),
                .input2(s_logisimNet34),
                .result(s_logisimNet195));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_26 (.input1(s_logisimNet27),
                .input2(s_logisimNet31),
                .result(s_logisimNet19));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_27 (.input1(s_logisimNet26),
                .input2(s_logisimNet3),
                .result(s_logisimNet60));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_28 (.input1(s_logisimNet307),
                .input2(s_logisimNet144),
                .result(s_logisimNet95));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_29 (.input1(s_logisimNet68),
                .input2(s_logisimNet273),
                .result(s_logisimNet256));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_30 (.input1(s_logisimNet227),
                .input2(s_logisimNet49),
                .result(s_logisimNet289));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_31 (.input1(s_logisimNet74),
                .input2(s_logisimNet64),
                .result(s_logisimNet140));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_32 (.input1(s_logisimNet140),
                .input2(s_logisimNet288),
                .result(s_logisimNet79));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_33 (.input1(s_logisimNet172),
                .input2(s_logisimNet168),
                .result(s_logisimNet320));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_34 (.input1(s_logisimNet197),
                .input2(s_logisimNet86),
                .result(s_logisimNet358));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_35 (.input1(s_logisimNet85),
                .input2(s_logisimNet3),
                .result(s_logisimNet318));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_36 (.input1(s_logisimNet4),
                .input2(s_logisimNet214),
                .result(s_logisimNet22));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_37 (.input1(s_logisimNet50),
                .input2(s_logisimNet102),
                .result(s_logisimNet374));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_38 (.input1(s_logisimNet299),
                .input2(s_logisimNet287),
                .result(s_logisimNet314));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_39 (.input1(s_logisimNet73),
                .input2(s_logisimNet46),
                .result(s_logisimNet82));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_40 (.input1(s_logisimNet74),
                .input2(s_logisimNet42),
                .result(s_logisimNet70));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_41 (.input1(s_logisimNet61),
                .input2(s_logisimNet15),
                .result(s_logisimNet306));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_42 (.input1(s_logisimNet50),
                .input2(s_logisimNet59),
                .result(s_logisimNet115));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_43 (.input1(s_logisimNet129),
                .input2(s_logisimNet202),
                .result(s_logisimNet307));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_44 (.input1(s_logisimNet14),
                .input2(s_logisimNet16),
                .result(s_logisimNet252));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_45 (.input1(s_logisimNet164),
                .input2(s_logisimNet317),
                .result(s_logisimNet353));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_46 (.input1(s_logisimNet17),
                .input2(s_logisimNet42),
                .result(s_logisimNet163));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_47 (.input1(s_logisimNet187),
                .input2(s_logisimNet314),
                .result(s_logisimNet110));

   Decoder_16   PLEXERS_48 (.decoderOut_0(s_logisimNet3),
                            .decoderOut_1(s_logisimNet29),
                            .decoderOut_10(s_logisimNet42),
                            .decoderOut_11(s_logisimNet7),
                            .decoderOut_12(s_logisimNet64),
                            .decoderOut_13(s_logisimNet32),
                            .decoderOut_14(s_logisimNet0),
                            .decoderOut_15(s_logisimNet59),
                            .decoderOut_2(s_logisimNet23),
                            .decoderOut_3(s_logisimNet46),
                            .decoderOut_4(s_logisimNet1),
                            .decoderOut_5(s_logisimNet31),
                            .decoderOut_6(s_logisimNet40),
                            .decoderOut_7(s_logisimNet102),
                            .decoderOut_8(s_logisimNet2),
                            .decoderOut_9(s_logisimNet15),
                            .enable(1'b1),
                            .sel(s_logisimBus100[7:4]));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_49 (.input1(s_logisimNet26),
                .input2(s_logisimNet1),
                .result(s_logisimNet202));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_50 (.input1(s_logisimNet175),
                .input2(s_logisimNet338),
                .result(s_logisimNet158));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_51 (.input1(s_logisimNet163),
                .input2(s_logisimNet9),
                .result(s_logisimNet47));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_52 (.input1(s_logisimNet4),
                .input2(s_logisimNet233),
                .result(s_logisimNet260));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_53 (.input1(s_logisimNet17),
                .input2(s_logisimNet1),
                .result(s_logisimNet186));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_54 (.input1(s_logisimNet74),
                .input2(s_logisimNet0),
                .result(s_logisimNet5));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_55 (.input1(s_logisimNet269),
                .input2(s_logisimNet351),
                .result(s_logisimNet89));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_56 (.input1(s_logisimNet75),
                .input2(s_logisimNet1),
                .result(s_logisimNet269));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_57 (.input1(s_logisimNet147),
                .input2(s_logisimNet194),
                .result(s_logisimNet148));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_58 (.input1(s_logisimNet146),
                .input2(s_logisimNet165),
                .result(s_logisimNet212));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_59 (.input1(s_logisimNet227),
                .input2(s_logisimNet117),
                .result(s_logisimNet276));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_60 (.input1(s_logisimNet96),
                .input2(s_logisimNet174),
                .result(s_logisimNet157));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_61 (.input1(s_logisimNet39),
                .input2(s_logisimNet286),
                .result(s_logisimNet119));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_62 (.input1(s_logisimNet27),
                .input2(s_logisimNet42),
                .result(s_logisimNet182));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_63 (.input1(s_logisimNet220),
                .input2(s_logisimNet60),
                .result(s_logisimNet284));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_64 (.input1(s_logisimNet167),
                .input2(s_logisimNet265),
                .result(s_logisimNet204));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_65 (.input1(s_logisimNet173),
                .input2(s_logisimNet297),
                .result(s_logisimNet126));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_66 (.input1(s_logisimNet67),
                .input2(s_logisimNet43),
                .result(s_logisimNet210));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_67 (.input1(s_logisimNet75),
                .input2(s_logisimNet29),
                .result(s_logisimNet328));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_68 (.input1(s_logisimNet73),
                .input2(s_logisimNet42),
                .result(s_logisimNet167));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_69 (.input1(s_logisimNet73),
                .input2(s_logisimNet102),
                .result(s_logisimNet35));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_70 (.input1(s_logisimNet138),
                .input2(s_logisimNet361),
                .result(s_logisimNet139));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_71 (.input1(s_logisimNet85),
                .input2(s_logisimNet1),
                .result(s_logisimNet238));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_72 (.input1(s_logisimNet75),
                .input2(s_logisimNet31),
                .result(s_logisimNet253));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_73 (.input1(s_logisimNet192),
                .input2(s_logisimNet345),
                .result(s_logisimNet159));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_74 (.input1(s_logisimNet181),
                .input2(s_logisimNet342),
                .result(s_logisimNet266));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_75 (.input1(s_logisimNet27),
                .input2(s_logisimNet0),
                .result(s_logisimNet236));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_76 (.input1(s_logisimNet149),
                .input2(s_logisimNet64),
                .result(s_logisimNet349));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_77 (.input1(s_logisimNet50),
                .input2(s_logisimNet1),
                .result(s_logisimNet66));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_78 (.input1(s_logisimNet10),
                .input2(s_logisimNet272),
                .result(s_logisimNet280));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_79 (.input1(s_logisimNet279),
                .input2(s_logisimNet263),
                .result(s_logisimNet317));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_80 (.input1(s_logisimNet50),
                .input2(s_logisimNet46),
                .result(s_logisimNet340));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_81 (.input1(s_logisimNet165),
                .input2(s_logisimNet336),
                .result(s_logisimNet351));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_82 (.input1(s_logisimNet53),
                .input2(s_logisimNet15),
                .result(s_logisimNet251));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_83 (.input1(s_logisimNet69),
                .input2(s_logisimNet281),
                .result(s_logisimNet310));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_84 (.input1(s_logisimNet87),
                .input2(s_logisimNet184),
                .result(s_logisimNet109));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_85 (.input1(s_logisimNet68),
                .input2(s_logisimNet241),
                .result(s_logisimNet45));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_86 (.input1(s_logisimNet208),
                .input2(s_logisimNet160),
                .result(s_logisimNet373));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_87 (.input1(s_logisimNet225),
                .input2(s_logisimNet192),
                .result(s_logisimNet274));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_88 (.input1(s_logisimNet26),
                .input2(s_logisimNet46),
                .result(s_logisimNet154));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_89 (.input1(s_logisimNet194),
                .input2(s_logisimNet333),
                .result(s_logisimNet155));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_90 (.input1(s_logisimNet20),
                .input2(s_logisimNet96),
                .result(s_logisimNet142));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_91 (.input1(s_logisimNet53),
                .input2(s_logisimNet42),
                .result(s_logisimNet13));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_92 (.input1(s_logisimNet243),
                .input2(s_logisimNet104),
                .result(s_logisimNet166));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_93 (.input1(s_logisimNet236),
                .input2(s_logisimNet157),
                .result(s_logisimNet350));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_94 (.input1(s_logisimNet234),
                .input2(s_logisimNet360),
                .result(s_logisimNet83));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_95 (.input1(s_logisimNet224),
                .input2(s_logisimNet275),
                .result(s_logisimNet332));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_96 (.input1(s_logisimNet162),
                .input2(s_logisimNet70),
                .result(s_logisimNet356));

   Decoder_16   PLEXERS_97 (.decoderOut_0(s_logisimNet73),
                            .decoderOut_1(s_logisimNet26),
                            .decoderOut_10(s_logisimNet149),
                            .decoderOut_11(),
                            .decoderOut_12(s_logisimNet74),
                            .decoderOut_13(s_logisimNet27),
                            .decoderOut_14(s_logisimNet17),
                            .decoderOut_15(),
                            .decoderOut_2(s_logisimNet313),
                            .decoderOut_3(),
                            .decoderOut_4(s_logisimNet61),
                            .decoderOut_5(s_logisimNet85),
                            .decoderOut_6(s_logisimNet53),
                            .decoderOut_7(),
                            .decoderOut_8(s_logisimNet50),
                            .decoderOut_9(s_logisimNet75),
                            .enable(1'b1),
                            .sel(s_logisimBus100[3:0]));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_98 (.input1(s_logisimNet318),
                .input2(s_logisimNet312),
                .result(s_logisimNet278));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_99 (.input1(s_logisimNet45),
                .input2(s_logisimNet230),
                .result(s_logisimNet78));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_100 (.input1(s_logisimNet260),
                 .input2(s_logisimNet358),
                 .result(s_logisimNet49));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_101 (.input1(s_logisimNet80),
                 .input2(s_logisimNet159),
                 .result(s_logisimNet247));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_102 (.input1(s_logisimNet143),
                 .input2(s_logisimNet164),
                 .result(s_logisimNet147));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_103 (.input1(s_logisimNet154),
                 .input2(s_logisimNet220),
                 .result(s_logisimNet245));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_104 (.input1(s_logisimNet27),
                 .input2(s_logisimNet64),
                 .result(s_logisimNet96));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_105 (.input1(s_logisimNet53),
                 .input2(s_logisimNet0),
                 .result(s_logisimNet218));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_106 (.input1(s_logisimNet75),
                 .input2(s_logisimNet32),
                 .result(s_logisimNet254));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_107 (.input1(s_logisimNet60),
                 .input2(s_logisimNet123),
                 .result(s_logisimNet24));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_108 (.input1(s_logisimNet90),
                 .input2(s_logisimNet296),
                 .result(s_logisimNet134));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_109 (.input1(s_logisimNet70),
                 .input2(s_logisimNet48),
                 .result(s_logisimNet288));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_110 (.input1(s_logisimNet84),
                 .input2(s_logisimNet122),
                 .result(s_logisimNet376));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_111 (.input1(s_logisimNet364),
                 .input2(s_logisimNet234),
                 .result(s_logisimNet348));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_112 (.input1(s_logisimNet73),
                 .input2(s_logisimNet3),
                 .result(s_logisimNet311));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_113 (.input1(s_logisimNet27),
                 .input2(s_logisimNet1),
                 .result(s_logisimNet170));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_114 (.input1(s_logisimNet213),
                 .input2(s_logisimNet361),
                 .result(s_logisimNet277));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_115 (.input1(s_logisimNet350),
                 .input2(s_logisimNet195),
                 .result(s_logisimNet343));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_116 (.input1(s_logisimNet104),
                 .input2(s_logisimNet334),
                 .result(s_logisimNet65));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_117 (.input1(s_logisimNet231),
                 .input2(s_logisimNet323),
                 .result(s_logisimNet272));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_118 (.input1(s_logisimNet182),
                 .input2(s_logisimNet315),
                 .result(s_logisimNet174));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_119 (.input1(s_logisimNet25),
                 .input2(s_logisimNet257),
                 .result(s_logisimNet237));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_120 (.input1(s_logisimNet50),
                 .input2(s_logisimNet42),
                 .result(s_logisimNet352));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_121 (.input1(s_logisimNet73),
                 .input2(s_logisimNet40),
                 .result(s_logisimNet380));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_122 (.input1(s_logisimNet53),
                 .input2(s_logisimNet2),
                 .result(s_logisimNet268));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_123 (.input1(s_logisimNet75),
                 .input2(s_logisimNet40),
                 .result(s_logisimNet56));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_124 (.input1(s_logisimNet53),
                 .input2(s_logisimNet3),
                 .result(s_logisimNet198));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_125 (.input1(s_logisimNet377),
                 .input2(s_logisimNet247),
                 .result(s_logisimNet322));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_126 (.input1(s_logisimNet39),
                 .input2(s_logisimNet236),
                 .result(s_logisimNet305));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_127 (.input1(s_logisimNet73),
                 .input2(s_logisimNet7),
                 .result(s_logisimNet188));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_128 (.input1(s_logisimNet149),
                 .input2(s_logisimNet1),
                 .result(s_logisimNet8));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_129 (.input1(s_logisimNet26),
                 .input2(s_logisimNet0),
                 .result(s_logisimNet179));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_130 (.input1(s_logisimNet130),
                 .input2(s_logisimNet304),
                 .result(s_logisimNet153));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_131 (.input1(s_logisimNet50),
                 .input2(s_logisimNet0),
                 .result(s_logisimNet262));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_132 (.input1(s_logisimNet53),
                 .input2(s_logisimNet7),
                 .result(s_logisimNet215));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_133 (.input1(s_logisimNet6),
                 .input2(s_logisimNet369),
                 .result(s_logisimNet189));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_134 (.input1(s_logisimNet128),
                 .input2(s_logisimNet47),
                 .result(s_logisimNet34));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_135 (.input1(s_logisimNet243),
                 .input2(s_logisimNet58),
                 .result(s_logisimNet214));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_136 (.input1(s_logisimNet232),
                 .input2(s_logisimNet150),
                 .result(s_logisimNet345));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_137 (.input1(s_logisimNet75),
                 .input2(s_logisimNet3),
                 .result(s_logisimNet336));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_138 (.input1(s_logisimNet50),
                 .input2(s_logisimNet32),
                 .result(s_logisimNet368));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_139 (.input1(s_logisimNet53),
                 .input2(s_logisimNet59),
                 .result(s_logisimNet239));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_140 (.input1(s_logisimNet209),
                 .input2(s_logisimNet131),
                 .result(s_logisimNet337));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_141 (.input1(s_logisimNet19),
                 .input2(s_logisimNet170),
                 .result(s_logisimNet141));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_142 (.input1(s_logisimNet85),
                 .input2(s_logisimNet42),
                 .result(s_logisimNet232));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_143 (.input1(s_logisimNet178),
                 .input2(s_logisimNet375),
                 .result(s_logisimNet325));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_144 (.input1(s_logisimNet50),
                 .input2(s_logisimNet3),
                 .result(s_logisimNet359));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_145 (.input1(s_logisimNet61),
                 .input2(s_logisimNet7),
                 .result(s_logisimNet205));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_146 (.input1(s_logisimNet26),
                 .input2(s_logisimNet2),
                 .result(s_logisimNet233));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_147 (.input1(s_logisimNet17),
                 .input2(s_logisimNet46),
                 .result(s_logisimNet113));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_148 (.input1(s_logisimNet8),
                 .input2(s_logisimNet283),
                 .result(s_logisimNet333));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_149 (.input1(s_logisimNet205),
                 .input2(s_logisimNet173),
                 .result(s_logisimNet265));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_150 (.input1(s_logisimNet73),
                 .input2(s_logisimNet15),
                 .result(s_logisimNet152));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_151 (.input1(s_logisimNet61),
                 .input2(s_logisimNet64),
                 .result(s_logisimNet97));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_152 (.input1(s_logisimNet253),
                 .input2(s_logisimNet269),
                 .result(s_logisimNet295));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_153 (.input1(s_logisimNet198),
                 .input2(s_logisimNet177),
                 .result(s_logisimNet319));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_154 (.input1(s_logisimNet17),
                 .input2(s_logisimNet3),
                 .result(s_logisimNet299));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_155 (.input1(s_logisimNet75),
                 .input2(s_logisimNet15),
                 .result(s_logisimNet227));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_156 (.input1(s_logisimNet99),
                 .input2(s_logisimNet135),
                 .result(s_logisimNet30));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_157 (.input1(s_logisimNet85),
                 .input2(s_logisimNet59),
                 .result(s_logisimNet181));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_158 (.input1(s_logisimNet97),
                 .input2(s_logisimNet126),
                 .result(s_logisimNet221));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_159 (.input1(s_logisimNet119),
                 .input2(s_logisimNet211),
                 .result(s_logisimNet200));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_160 (.input1(s_logisimNet50),
                 .input2(s_logisimNet40),
                 .result(s_logisimNet219));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_161 (.input1(s_logisimNet61),
                 .input2(s_logisimNet42),
                 .result(s_logisimNet173));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_162 (.input1(s_logisimNet16),
                 .input2(s_logisimNet12),
                 .result(s_logisimNet196));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_163 (.input1(s_logisimNet26),
                 .input2(s_logisimNet40),
                 .result(s_logisimNet104));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_164 (.input1(s_logisimNet134),
                 .input2(s_logisimNet142),
                 .result(s_logisimNet330));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_165 (.input1(s_logisimNet53),
                 .input2(s_logisimNet40),
                 .result(s_logisimNet164));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_166 (.input1(s_logisimNet50),
                 .input2(s_logisimNet31),
                 .result(s_logisimNet367));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_167 (.input1(s_logisimNet95),
                 .input2(s_logisimNet295),
                 .result(s_logisimNet133));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_168 (.input1(s_logisimNet188),
                 .input2(s_logisimNet217),
                 .result(s_logisimNet190));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_169 (.input1(s_logisimNet149),
                 .input2(s_logisimNet2),
                 .result(s_logisimNet62));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_170 (.input1(s_logisimNet50),
                 .input2(s_logisimNet15),
                 .result(s_logisimNet127));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_171 (.input1(s_logisimNet172),
                 .input2(s_logisimNet128),
                 .result(s_logisimNet230));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_172 (.input1(s_logisimNet85),
                 .input2(s_logisimNet29),
                 .result(s_logisimNet312));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_173 (.input1(s_logisimNet84),
                 .input2(s_logisimNet312),
                 .result(s_logisimNet275));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_174 (.input1(s_logisimNet113),
                 .input2(s_logisimNet290),
                 .result(s_logisimNet92));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_175 (.input1(s_logisimNet120),
                 .input2(s_logisimNet93),
                 .result(s_logisimNet339));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_176 (.input1(s_logisimNet130),
                 .input2(s_logisimNet271),
                 .result(s_logisimNet183));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_177 (.input1(s_logisimNet216),
                 .input2(s_logisimNet36),
                 .result(s_logisimNet285));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_178 (.input1(s_logisimNet75),
                 .input2(s_logisimNet42),
                 .result(s_logisimNet255));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_179 (.input1(s_logisimNet27),
                 .input2(s_logisimNet46),
                 .result(s_logisimNet138));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_180 (.input1(s_logisimNet105),
                 .input2(s_logisimNet249),
                 .result(s_logisimNet309));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_181 (.input1(s_logisimNet204),
                 .input2(s_logisimNet356),
                 .result(s_logisimNet124));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_182 (.input1(s_logisimNet75),
                 .input2(s_logisimNet23),
                 .result(s_logisimNet165));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_183 (.input1(s_logisimNet143),
                 .input2(s_logisimNet210),
                 .result(s_logisimNet292));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_184 (.input1(s_logisimNet166),
                 .input2(s_logisimNet252),
                 .result(s_logisimNet175));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_185 (.input1(s_logisimNet149),
                 .input2(s_logisimNet40),
                 .result(s_logisimNet194));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_186 (.input1(s_logisimNet27),
                 .input2(s_logisimNet32),
                 .result(s_logisimNet20));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_187 (.input1(s_logisimNet131),
                 .input2(s_logisimNet132),
                 .result(s_logisimNet9));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_188 (.input1(s_logisimNet348),
                 .input2(s_logisimNet280),
                 .result(s_logisimNet371));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_189 (.input1(s_logisimNet69),
                 .input2(s_logisimNet309),
                 .result(s_logisimNet116));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_190 (.input1(s_logisimNet75),
                 .input2(s_logisimNet64),
                 .result(s_logisimNet231));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_191 (.input1(s_logisimNet85),
                 .input2(s_logisimNet46),
                 .result(s_logisimNet84));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_192 (.input1(s_logisimNet238),
                 .input2(s_logisimNet344),
                 .result(s_logisimNet12));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_193 (.input1(s_logisimNet118),
                 .input2(s_logisimNet167),
                 .result(s_logisimNet264));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_194 (.input1(s_logisimNet105),
                 .input2(s_logisimNet185),
                 .result(s_logisimNet250));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_195 (.input1(s_logisimNet26),
                 .input2(s_logisimNet32),
                 .result(s_logisimNet130));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_196 (.input1(s_logisimNet222),
                 .input2(s_logisimNet108),
                 .result(s_logisimNet235));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_197 (.input1(s_logisimNet61),
                 .input2(s_logisimNet0),
                 .result(s_logisimNet203));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_198 (.input1(s_logisimNet27),
                 .input2(s_logisimNet3),
                 .result(s_logisimNet213));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_199 (.input1(s_logisimNet297),
                 .input2(s_logisimNet306),
                 .result(s_logisimNet99));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_200 (.input1(s_logisimNet270),
                 .input2(s_logisimNet300),
                 .result(s_logisimNet168));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_201 (.input1(s_logisimNet14),
                 .input2(s_logisimNet332),
                 .result(s_logisimNet52));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_202 (.input1(s_logisimNet20),
                 .input2(s_logisimNet38),
                 .result(s_logisimNet286));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_203 (.input1(s_logisimNet44),
                 .input2(s_logisimNet8),
                 .result(s_logisimNet111));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_204 (.input1(s_logisimNet181),
                 .input2(s_logisimNet80),
                 .result(s_logisimNet355));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_205 (.input1(s_logisimNet183),
                 .input2(s_logisimNet274),
                 .result(s_logisimNet90));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_206 (.input1(s_logisimNet87),
                 .input2(s_logisimNet177),
                 .result(s_logisimNet43));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_207 (.input1(s_logisimNet50),
                 .input2(s_logisimNet23),
                 .result(s_logisimNet372));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_208 (.input1(s_logisimNet54),
                 .input2(s_logisimNet246),
                 .result(s_logisimNet283));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_209 (.input1(s_logisimNet27),
                 .input2(s_logisimNet40),
                 .result(s_logisimNet185));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_210 (.input1(s_logisimNet27),
                 .input2(s_logisimNet15),
                 .result(s_logisimNet69));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_211 (.input1(s_logisimNet251),
                 .input2(s_logisimNet268),
                 .result(s_logisimNet209));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_212 (.input1(s_logisimNet242),
                 .input2(s_logisimNet339),
                 .result(s_logisimNet180));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_213 (.input1(s_logisimNet225),
                 .input2(s_logisimNet237),
                 .result(s_logisimNet342));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_214 (.input1(s_logisimNet73),
                 .input2(s_logisimNet23),
                 .result(s_logisimNet160));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_215 (.input1(s_logisimNet254),
                 .input2(s_logisimNet231),
                 .result(s_logisimNet296));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_216 (.input1(s_logisimNet67),
                 .input2(s_logisimNet279),
                 .result(s_logisimNet44));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_217 (.input1(s_logisimNet149),
                 .input2(s_logisimNet23),
                 .result(s_logisimNet54));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_218 (.input1(s_logisimNet85),
                 .input2(s_logisimNet32),
                 .result(s_logisimNet225));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_219 (.input1(s_logisimNet26),
                 .input2(s_logisimNet23),
                 .result(s_logisimNet220));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_220 (.input1(s_logisimNet253),
                 .input2(s_logisimNet291),
                 .result(s_logisimNet21));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_221 (.input1(s_logisimNet17),
                 .input2(s_logisimNet64),
                 .result(s_logisimNet128));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_222 (.input1(s_logisimNet241),
                 .input2(s_logisimNet169),
                 .result(s_logisimNet316));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_223 (.input1(s_logisimNet50),
                 .input2(s_logisimNet2),
                 .result(s_logisimNet298));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_224 (.input1(s_logisimNet61),
                 .input2(s_logisimNet2),
                 .result(s_logisimNet297));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_225 (.input1(s_logisimNet106),
                 .input2(s_logisimNet22),
                 .result(s_logisimNet304));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_226 (.input1(s_logisimNet138),
                 .input2(s_logisimNet33),
                 .result(s_logisimNet375));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_227 (.input1(s_logisimNet186),
                 .input2(s_logisimNet326),
                 .result(s_logisimNet57));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_228 (.input1(s_logisimNet71),
                 .input2(s_logisimNet212),
                 .result(s_logisimNet178));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_229 (.input1(s_logisimNet27),
                 .input2(s_logisimNet59),
                 .result(s_logisimNet39));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_230 (.input1(s_logisimNet216),
                 .input2(s_logisimNet10),
                 .result(s_logisimNet362));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_231 (.input1(s_logisimNet91),
                 .input2(s_logisimNet21),
                 .result(s_logisimNet117));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_232 (.input1(s_logisimNet73),
                 .input2(s_logisimNet32),
                 .result(s_logisimNet223));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_233 (.input1(s_logisimNet73),
                 .input2(s_logisimNet64),
                 .result(s_logisimNet118));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_234 (.input1(s_logisimNet50),
                 .input2(s_logisimNet7),
                 .result(s_logisimNet303));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_235 (.input1(s_logisimNet26),
                 .input2(s_logisimNet7),
                 .result(s_logisimNet106));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_236 (.input1(s_logisimNet207),
                 .input2(s_logisimNet176),
                 .result(s_logisimNet382));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_237 (.input1(s_logisimNet73),
                 .input2(s_logisimNet59),
                 .result(s_logisimNet137));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_238 (.input1(s_logisimNet129),
                 .input2(s_logisimNet329),
                 .result(s_logisimNet58));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_239 (.input1(s_logisimNet98),
                 .input2(s_logisimNet276),
                 .result(s_logisimNet261));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_240 (.input1(s_logisimNet171),
                 .input2(s_logisimNet228),
                 .result(s_logisimNet300));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_241 (.input1(s_logisimNet122),
                 .input2(s_logisimNet318),
                 .result(s_logisimNet344));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_242 (.input1(s_logisimNet373),
                 .input2(s_logisimNet343),
                 .result(s_logisimNet354));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_243 (.input1(s_logisimNet244),
                 .input2(s_logisimNet140),
                 .result(s_logisimNet294));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_244 (.input1(s_logisimNet53),
                 .input2(s_logisimNet102),
                 .result(s_logisimNet143));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_245 (.input1(s_logisimNet170),
                 .input2(s_logisimNet206),
                 .result(s_logisimNet156));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_246 (.input1(s_logisimNet17),
                 .input2(s_logisimNet32),
                 .result(s_logisimNet172));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_247 (.input1(s_logisimNet77),
                 .input2(s_logisimNet264),
                 .result(s_logisimNet364));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_248 (.input1(s_logisimNet85),
                 .input2(s_logisimNet31),
                 .result(s_logisimNet224));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_249 (.input1(s_logisimNet25),
                 .input2(s_logisimNet232),
                 .result(s_logisimNet381));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_250 (.input1(s_logisimNet41),
                 .input2(s_logisimNet179),
                 .result(s_logisimNet248));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_251 (.input1(s_logisimNet26),
                 .input2(s_logisimNet15),
                 .result(s_logisimNet4));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_252 (.input1(s_logisimNet293),
                 .input2(s_logisimNet116),
                 .result(s_logisimNet38));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_253 (.input1(s_logisimNet152),
                 .input2(s_logisimNet101),
                 .result(s_logisimNet217));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_254 (.input1(s_logisimNet193),
                 .input2(s_logisimNet92),
                 .result(s_logisimNet191));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_255 (.input1(s_logisimNet75),
                 .input2(s_logisimNet59),
                 .result(s_logisimNet216));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_256 (.input1(s_logisimNet75),
                 .input2(s_logisimNet7),
                 .result(s_logisimNet98));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_257 (.input1(s_logisimNet50),
                 .input2(s_logisimNet64),
                 .result(s_logisimNet379));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_258 (.input1(s_logisimNet223),
                 .input2(s_logisimNet190),
                 .result(s_logisimNet331));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_259 (.input1(s_logisimNet85),
                 .input2(s_logisimNet102),
                 .result(s_logisimNet14));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_260 (.input1(s_logisimNet114),
                 .input2(s_logisimNet266),
                 .result(s_logisimNet366));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_261 (.input1(s_logisimNet75),
                 .input2(s_logisimNet102),
                 .result(s_logisimNet91));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_262 (.input1(s_logisimNet26),
                 .input2(s_logisimNet31),
                 .result(s_logisimNet129));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_263 (.input1(s_logisimNet74),
                 .input2(s_logisimNet7),
                 .result(s_logisimNet162));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_264 (.input1(s_logisimNet251),
                 .input2(s_logisimNet292),
                 .result(s_logisimNet37));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_265 (.input1(s_logisimNet179),
                 .input2(s_logisimNet335),
                 .result(s_logisimNet378));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_266 (.input1(s_logisimNet254),
                 .input2(s_logisimNet261),
                 .result(s_logisimNet36));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_267 (.input1(s_logisimNet26),
                 .input2(s_logisimNet59),
                 .result(s_logisimNet41));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_268 (.input1(s_logisimNet85),
                 .input2(s_logisimNet23),
                 .result(s_logisimNet122));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_269 (.input1(s_logisimNet203),
                 .input2(s_logisimNet221),
                 .result(s_logisimNet341));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_270 (.input1(s_logisimNet73),
                 .input2(s_logisimNet1),
                 .result(s_logisimNet370));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_271 (.input1(s_logisimNet149),
                 .input2(s_logisimNet15),
                 .result(s_logisimNet365));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_272 (.input1(s_logisimNet199),
                 .input2(s_logisimNet277),
                 .result(s_logisimNet121));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_273 (.input1(s_logisimNet336),
                 .input2(s_logisimNet328),
                 .result(s_logisimNet347));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_274 (.input1(s_logisimNet17),
                 .input2(s_logisimNet23),
                 .result(s_logisimNet290));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_275 (.input1(s_logisimNet53),
                 .input2(s_logisimNet23),
                 .result(s_logisimNet184));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_276 (.input1(s_logisimNet109),
                 .input2(s_logisimNet54),
                 .result(s_logisimNet193));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_277 (.input1(s_logisimNet24),
                 .input2(s_logisimNet278),
                 .result(s_logisimNet18));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_278 (.input1(s_logisimNet245),
                 .input2(s_logisimNet376),
                 .result(s_logisimNet71));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_279 (.input1(s_logisimNet75),
                 .input2(s_logisimNet46),
                 .result(s_logisimNet146));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_280 (.input1(s_logisimNet53),
                 .input2(s_logisimNet1),
                 .result(s_logisimNet279));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_281 (.input1(s_logisimNet18),
                 .input2(s_logisimNet347),
                 .result(s_logisimNet199));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_282 (.input1(s_logisimNet26),
                 .input2(s_logisimNet102),
                 .result(s_logisimNet243));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_283 (.input1(s_logisimNet171),
                 .input2(s_logisimNet186),
                 .result(s_logisimNet229));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_284 (.input1(s_logisimNet53),
                 .input2(s_logisimNet46),
                 .result(s_logisimNet87));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_285 (.input1(s_logisimNet233),
                 .input2(s_logisimNet65),
                 .result(s_logisimNet145));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_286 (.input1(s_logisimNet13),
                 .input2(s_logisimNet88),
                 .result(s_logisimNet169));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_287 (.input1(s_logisimNet268),
                 .input2(s_logisimNet353),
                 .result(s_logisimNet88));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_288 (.input1(s_logisimNet98),
                 .input2(s_logisimNet255),
                 .result(s_logisimNet72));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_289 (.input1(s_logisimNet197),
                 .input2(s_logisimNet52),
                 .result(s_logisimNet257));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_290 (.input1(s_logisimNet17),
                 .input2(s_logisimNet40),
                 .result(s_logisimNet282));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_291 (.input1(s_logisimNet282),
                 .input2(s_logisimNet57),
                 .result(s_logisimNet132));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_292 (.input1(s_logisimNet215),
                 .input2(s_logisimNet13),
                 .result(s_logisimNet360));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_293 (.input1(s_logisimNet85),
                 .input2(s_logisimNet15),
                 .result(s_logisimNet197));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_294 (.input1(s_logisimNet91),
                 .input2(s_logisimNet56),
                 .result(s_logisimNet338));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_295 (.input1(s_logisimNet19),
                 .input2(s_logisimNet139),
                 .result(s_logisimNet249));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_296 (.input1(s_logisimNet17),
                 .input2(s_logisimNet59),
                 .result(s_logisimNet120));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_297 (.input1(s_logisimNet158),
                 .input2(s_logisimNet250),
                 .result(s_logisimNet28));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_298 (.input1(s_logisimNet74),
                 .input2(s_logisimNet40),
                 .result(s_logisimNet176));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_299 (.input1(s_logisimNet203),
                 .input2(s_logisimNet77),
                 .result(s_logisimNet151));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_300 (.input1(s_logisimNet50),
                 .input2(s_logisimNet29),
                 .result(s_logisimNet302));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_301 (.input1(s_logisimNet239),
                 .input2(s_logisimNet256),
                 .result(s_logisimNet114));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_302 (.input1(s_logisimNet73),
                 .input2(s_logisimNet29),
                 .result(s_logisimNet51));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_303 (.input1(s_logisimNet281),
                 .input2(s_logisimNet259),
                 .result(s_logisimNet315));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_304 (.input1(s_logisimNet17),
                 .input2(s_logisimNet31),
                 .result(s_logisimNet171));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_305 (.input1(s_logisimNet53),
                 .input2(s_logisimNet31),
                 .result(s_logisimNet67));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_306 (.input1(s_logisimNet26),
                 .input2(s_logisimNet29),
                 .result(s_logisimNet123));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_307 (.input1(s_logisimNet137),
                 .input2(s_logisimNet331),
                 .result(s_logisimNet267));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_308 (.input1(s_logisimNet26),
                 .input2(s_logisimNet42),
                 .result(s_logisimNet81));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_309 (.input1(s_logisimNet215),
                 .input2(s_logisimNet37),
                 .result(s_logisimNet273));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_310 (.input1(s_logisimNet74),
                 .input2(s_logisimNet2),
                 .result(s_logisimNet135));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_311 (.input1(s_logisimNet146),
                 .input2(s_logisimNet328),
                 .result(s_logisimNet291));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_312 (.input1(s_logisimNet55),
                 .input2(s_logisimNet381),
                 .result(s_logisimNet346));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_313 (.input1(s_logisimNet184),
                 .input2(s_logisimNet198),
                 .result(s_logisimNet263));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_314 (.input1(s_logisimNet154),
                 .input2(s_logisimNet123),
                 .result(s_logisimNet329));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_315 (.input1(s_logisimNet319),
                 .input2(s_logisimNet246),
                 .result(s_logisimNet187));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_316 (.input1(s_logisimNet17),
                 .input2(s_logisimNet2),
                 .result(s_logisimNet131));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_317 (.input1(s_logisimNet293),
                 .input2(s_logisimNet182),
                 .result(s_logisimNet369));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_318 (.input1(s_logisimNet27),
                 .input2(s_logisimNet7),
                 .result(s_logisimNet293));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_319 (.input1(s_logisimNet205),
                 .input2(s_logisimNet306),
                 .result(s_logisimNet107));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_320 (.input1(s_logisimNet53),
                 .input2(s_logisimNet29),
                 .result(s_logisimNet177));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_321 (.input1(s_logisimNet248),
                 .input2(s_logisimNet355),
                 .result(s_logisimNet240));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_322 (.input1(s_logisimNet86),
                 .input2(s_logisimNet196),
                 .result(s_logisimNet150));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_323 (.input1(s_logisimNet161),
                 .input2(s_logisimNet163),
                 .result(s_logisimNet321));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_324 (.input1(s_logisimNet85),
                 .input2(s_logisimNet2),
                 .result(s_logisimNet86));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_325 (.input1(s_logisimNet240),
                 .input2(s_logisimNet362),
                 .result(s_logisimNet103));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_326 (.input1(s_logisimNet289),
                 .input2(s_logisimNet310),
                 .result(s_logisimNet327));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_327 (.input1(s_logisimNet53),
                 .input2(s_logisimNet64),
                 .result(s_logisimNet241));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_328 (.input1(s_logisimNet135),
                 .input2(s_logisimNet207),
                 .result(s_logisimNet48));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_329 (.input1(s_logisimNet133),
                 .input2(s_logisimNet141),
                 .result(s_logisimNet357));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_330 (.input1(s_logisimNet271),
                 .input2(s_logisimNet201),
                 .result(s_logisimNet335));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_331 (.input1(s_logisimNet83),
                 .input2(s_logisimNet321),
                 .result(s_logisimNet125));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_332 (.input1(s_logisimNet346),
                 .input2(s_logisimNet72),
                 .result(s_logisimNet6));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_333 (.input1(s_logisimNet239),
                 .input2(s_logisimNet218),
                 .result(s_logisimNet242));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_334 (.input1(s_logisimNet81),
                 .input2(s_logisimNet145),
                 .result(s_logisimNet201));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_335 (.input1(s_logisimNet149),
                 .input2(s_logisimNet3),
                 .result(s_logisimNet246));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_336 (.input1(s_logisimNet120),
                 .input2(s_logisimNet320),
                 .result(s_logisimNet211));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_337 (.input1(s_logisimNet224),
                 .input2(s_logisimNet238),
                 .result(s_logisimNet144));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_338 (.input1(1'b0),
                 .input2(s_logisimNet284),
                 .result(s_logisimNet334));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_339 (.input1(s_logisimNet73),
                 .input2(s_logisimNet0),
                 .result(s_logisimNet77));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_340 (.input1(s_logisimNet17),
                 .input2(s_logisimNet29),
                 .result(s_logisimNet287));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_341 (.input1(s_logisimNet27),
                 .input2(s_logisimNet2),
                 .result(s_logisimNet281));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_342 (.input1(s_logisimNet148),
                 .input2(s_logisimNet301),
                 .result(s_logisimNet11));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_343 (.input1(s_logisimNet149),
                 .input2(s_logisimNet42),
                 .result(s_logisimNet258));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_344 (.input1(s_logisimNet5),
                 .input2(s_logisimNet79),
                 .result(s_logisimNet208));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_345 (.input1(s_logisimNet85),
                 .input2(s_logisimNet40),
                 .result(s_logisimNet16));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_346 (.input1(s_logisimNet17),
                 .input2(s_logisimNet102),
                 .result(s_logisimNet270));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_347 (.input1(s_logisimNet73),
                 .input2(s_logisimNet31),
                 .result(s_logisimNet222));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_348 (.input1(s_logisimNet185),
                 .input2(s_logisimNet156),
                 .result(s_logisimNet259));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_349 (.input1(s_logisimNet270),
                 .input2(s_logisimNet282),
                 .result(s_logisimNet301));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_350 (.input1(s_logisimNet41),
                 .input2(s_logisimNet153),
                 .result(s_logisimNet324));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_351 (.input1(s_logisimNet17),
                 .input2(s_logisimNet7),
                 .result(s_logisimNet161));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_352 (.input1(s_logisimNet107),
                 .input2(s_logisimNet366),
                 .result(s_logisimNet363));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_353 (.input1(s_logisimNet27),
                 .input2(s_logisimNet23),
                 .result(s_logisimNet33));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_354 (.input1(s_logisimNet341),
                 .input2(s_logisimNet322),
                 .result(s_logisimNet308));


endmodule
