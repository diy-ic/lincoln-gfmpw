magic
tech gf180mcuD
magscale 1 5
timestamp 1702054272
<< obsm1 >>
rect 672 1538 57960 58830
<< metal2 >>
rect 27552 0 27608 400
rect 27888 0 27944 400
rect 30576 0 30632 400
rect 35280 0 35336 400
<< obsm2 >>
rect 966 430 57778 58819
rect 966 400 27522 430
rect 27638 400 27858 430
rect 27974 400 30546 430
rect 30662 400 35250 430
rect 35366 400 57778 430
<< metal3 >>
rect 0 56112 400 56168
<< obsm3 >>
rect 400 56198 57783 58814
rect 430 56082 57783 56198
rect 400 1554 57783 56082
<< metal4 >>
rect 2224 1538 2384 58830
rect 9904 1538 10064 58830
rect 17584 1538 17744 58830
rect 25264 1538 25424 58830
rect 32944 1538 33104 58830
rect 40624 1538 40784 58830
rect 48304 1538 48464 58830
rect 55984 1538 56144 58830
<< obsm4 >>
rect 1526 3369 2194 57279
rect 2414 3369 9874 57279
rect 10094 3369 17554 57279
rect 17774 3369 25234 57279
rect 25454 3369 32914 57279
rect 33134 3369 40594 57279
rect 40814 3369 48274 57279
rect 48494 3369 54474 57279
<< labels >>
rlabel metal2 s 27552 0 27608 400 6 spi_clock_i
port 1 nsew signal input
rlabel metal2 s 27888 0 27944 400 6 spi_cs_i
port 2 nsew signal input
rlabel metal2 s 35280 0 35336 400 6 spi_pico_i
port 3 nsew signal input
rlabel metal2 s 30576 0 30632 400 6 spi_poci_o
port 4 nsew signal output
rlabel metal3 s 0 56112 400 56168 6 sys_clock_i
port 5 nsew signal input
rlabel metal4 s 2224 1538 2384 58830 6 vdd
port 6 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58830 6 vdd
port 6 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58830 6 vdd
port 6 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58830 6 vdd
port 6 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58830 6 vss
port 7 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58830 6 vss
port 7 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58830 6 vss
port 7 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58830 6 vss
port 7 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 58680 60472
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9706600
string GDS_FILE /home/kris/repos/diy-ic/lincoln-gfmpw-1d/openlane/titan/runs/23_12_08_16_45/results/signoff/titan.magic.gds
string GDS_START 455504
<< end >>

