magic
tech gf180mcuD
magscale 1 5
timestamp 1701617586
<< obsm1 >>
rect 672 1538 50680 51382
<< metal2 >>
rect 26880 0 26936 400
rect 34944 0 35000 400
rect 36624 0 36680 400
rect 38304 0 38360 400
<< obsm2 >>
rect 686 430 50610 51371
rect 686 400 26850 430
rect 26966 400 34914 430
rect 35030 400 36594 430
rect 36710 400 38274 430
rect 38390 400 50610 430
<< metal3 >>
rect 0 50736 400 50792
<< obsm3 >>
rect 400 50822 50559 51366
rect 430 50706 50559 50822
rect 400 1554 50559 50706
<< metal4 >>
rect 2224 1538 2384 51382
rect 9904 1538 10064 51382
rect 17584 1538 17744 51382
rect 25264 1538 25424 51382
rect 32944 1538 33104 51382
rect 40624 1538 40784 51382
rect 48304 1538 48464 51382
<< obsm4 >>
rect 4998 2417 9874 50839
rect 10094 2417 17554 50839
rect 17774 2417 25234 50839
rect 25454 2417 32914 50839
rect 33134 2417 40594 50839
rect 40814 2417 47138 50839
<< labels >>
rlabel metal2 s 34944 0 35000 400 6 spi_clock_i
port 1 nsew signal input
rlabel metal2 s 36624 0 36680 400 6 spi_cs_i
port 2 nsew signal input
rlabel metal2 s 26880 0 26936 400 6 spi_pico_i
port 3 nsew signal input
rlabel metal2 s 38304 0 38360 400 6 spi_poci_o
port 4 nsew signal output
rlabel metal3 s 0 50736 400 50792 6 sys_clock_i
port 5 nsew signal input
rlabel metal4 s 2224 1538 2384 51382 6 vdd
port 6 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 51382 6 vdd
port 6 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 51382 6 vdd
port 6 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 51382 6 vdd
port 6 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 51382 6 vss
port 7 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 51382 6 vss
port 7 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 51382 6 vss
port 7 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 51369 53161
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8669832
string GDS_FILE /home/kris/repos/diy-ic/lincoln-gfmpw/openlane/titan/runs/23_12_03_15_28/results/signoff/titan.magic.gds
string GDS_START 474308
<< end >>

