* NGSPICE file created from titan.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

.subckt titan spi_clock_i spi_cs_i spi_pico_i spi_poci_o sys_clock_i vdd vss
X_05903_ _01561_ _01562_ _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06883_ _02418_ _02461_ _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_126_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09671_ _00258_ net260 ci_neuron.uut_simple_neuron.x3\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05834_ _01162_ _01200_ _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout56_I net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08622_ _03889_ _03879_ _04081_ _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05765_ _01427_ _01428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_25_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08553_ ci_neuron.value_i\[15\] _04001_ _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07504_ _03123_ _03130_ _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_85_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08484_ _03968_ _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07435_ _02979_ _03060_ _03062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05696_ _01252_ _01324_ _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07366_ _02962_ _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07297_ _02873_ _02877_ _02925_ _02926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06317_ ci_neuron.uut_simple_neuron.x3\[8\] _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09105_ _04360_ _04445_ _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06248_ _01877_ _01896_ _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05076__A2 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09036_ _04361_ _04383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06179_ _01827_ _01830_ _01831_ _01832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_102_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09211__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09938_ _00453_ net168 ci_neuron.uut_simple_neuron.x0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09869_ _00060_ net33 ci_neuron.value_i\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09373__S1 _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09202__A1 _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10009_ ci_neuron.input_memory\[1\]\[9\] net205 ci_neuron.uut_simple_neuron.titan_id_1\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05550_ _00859_ _01178_ _01174_ _01218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_121_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05451__I _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05481_ _01097_ _01150_ _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07220_ _02789_ _02848_ _02849_ _02850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08619__I1 _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07151_ _02718_ _02759_ _02782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06102_ _00747_ ci_neuron.uut_simple_neuron.x2\[29\] _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09441__A1 ci_neuron.output_memory\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07082_ _01835_ _02713_ _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06033_ _01650_ _01679_ _01690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout116 net117 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout127 net135 net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout138 net140 net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout105 net106 net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout149 net150 net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07984_ ci_neuron.uut_simple_neuron.titan_id_2\[26\] ci_neuron.uut_simple_neuron.titan_id_5\[26\]
+ _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_38_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06935_ _02472_ _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08555__I0 _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09723_ _00302_ net256 ci_neuron.uut_simple_neuron.x2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_2_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06866_ _02388_ _02501_ _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_87_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09654_ _04810_ _04826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05817_ _01327_ _01478_ _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08605_ _03864_ _04077_ _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06797_ _02376_ _02432_ _02433_ _02434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09585_ _04607_ ci_neuron.normalised_stream_write_address\[1\] _04785_ _04787_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05748_ _01361_ _01409_ _01410_ _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08536_ _04024_ _00262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05679_ _01342_ _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08467_ _03950_ _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08483__A2 _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07418_ _01988_ _01991_ _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08398_ _03902_ _00188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07349_ _02974_ _02977_ _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_98_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09283__I1 ci_neuron.input_memory\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09019_ internal_ih.data_pointer\[1\] _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09499__A1 ci_neuron.output_memory\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04980__A1 internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_107_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06237__A1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06788__A2 _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05212__A2 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04981_ _00684_ _00039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06720_ _02358_ _00235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08757__I _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04971__A1 internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06651_ _02044_ _02290_ _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05602_ _00937_ _01266_ _01268_ _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_69_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06582_ _02188_ _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05181__I _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09370_ _04604_ _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_35_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05533_ _01123_ _01162_ _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_82_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08321_ ci_neuron.uut_simple_neuron.x0\[18\] _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05464_ _01131_ _01107_ _01133_ _01056_ _01134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_08252_ _03775_ _00199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_15_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07203_ _02784_ _02833_ _02834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_6_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05395_ _00934_ _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08183_ _03692_ _03700_ _03712_ _03716_ _03717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_40_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07134_ _02647_ _02765_ _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07065_ _02652_ _02697_ _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06016_ _01665_ _01673_ _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09568__I2 _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07967_ _03537_ _00142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06918_ _02498_ _02552_ _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08528__I0 _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09706_ _00285_ net131 internal_ih.spi_rx_byte_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07898_ ci_neuron.uut_simple_neuron.titan_id_2\[11\] ci_neuron.uut_simple_neuron.titan_id_5\[11\]
+ _03480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04962__A1 internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06703__A2 _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06849_ _02440_ _02456_ _02485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09637_ ci_neuron.stream_o\[20\] ci_neuron.output_memory\[20\] _04816_ _04817_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09568_ _03915_ ci_neuron.input_memory\[1\]\[29\] _01751_ ci_neuron.uut_simple_neuron.x3\[29\]
+ _04760_ _04761_ _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_38_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08519_ ci_neuron.value_i\[10\] _03971_ _04009_ _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_93_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09499_ ci_neuron.output_memory\[19\] _04698_ _04715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09405__A1 ci_neuron.output_memory\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09256__I1 ci_neuron.uut_simple_neuron.x0\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06219__A1 _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10274_ _00567_ net142 ci_neuron.stream_o\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_14_Left_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_12_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05180_ net38 _00837_ _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08870_ _04276_ _00344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07821_ ci_neuron.uut_simple_neuron.titan_id_4\[30\] ci_neuron.uut_simple_neuron.titan_id_3\[30\]
+ _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07752_ ci_neuron.uut_simple_neuron.titan_id_4\[18\] ci_neuron.uut_simple_neuron.titan_id_3\[18\]
+ _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04964_ _00664_ _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06703_ _02332_ _02341_ _02342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_79_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07683_ _03301_ _00123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04895_ _00627_ _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06634_ _01907_ _02273_ _02274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06697__A1 _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08930__I0 internal_ih.byte5\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09422_ _04597_ _04649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09353_ internal_ih.expected_byte_count\[3\] _04352_ _04590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06565_ _02203_ _02206_ _02207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06449__A1 _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08304_ _03820_ _00176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06496_ _02094_ _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05516_ _01096_ _01149_ _01184_ _01185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09284_ _04551_ _00483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05447_ _01116_ _01117_ _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08235_ _03752_ ci_neuron.uut_simple_neuron.x0\[7\] _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_15_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05378_ _01012_ _01020_ _00961_ _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08166_ _03696_ _03701_ _03702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07117_ _02175_ _02193_ _02749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08097_ _03643_ _03645_ _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07048_ ci_neuron.uut_simple_neuron.x3\[21\] ci_neuron.uut_simple_neuron.x3\[22\]
+ _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08999_ internal_ih.current_instruction\[7\] _04341_ _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_98_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_50_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08601__A2 _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10257_ _00000_ net68 ci_neuron.stream_enabled vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10188_ _00086_ net44 ci_neuron.uut_simple_neuron.titan_id_2\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08912__I0 internal_ih.byte4\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07340__A2 _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06350_ _01994_ _01995_ _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_127_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06281_ _01928_ _01929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05301_ ci_neuron.uut_simple_neuron.x2\[7\] ci_neuron.uut_simple_neuron.x2\[8\] _00975_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05232_ _00894_ _00897_ _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08770__I _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08020_ ci_neuron.uut_simple_neuron.titan_id_1\[3\] ci_neuron.uut_simple_neuron.titan_id_0\[3\]
+ _03580_ _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_102_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05163_ _00840_ _00841_ _00842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_4_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout7 net8 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05094_ _00736_ _00774_ _00775_ _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09971_ _00486_ net179 ci_neuron.input_memory\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08922_ _04305_ _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_90_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08853_ _04266_ _00337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07804_ _03399_ _03401_ _03402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_98_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05996_ _01609_ _01627_ _01653_ _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08784_ _00911_ _04221_ _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04917__B2 internal_ih.byte1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07735_ _03344_ _00102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05590__A1 _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04947_ internal_ih.byte0\[0\] _00665_ _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08903__I0 internal_ih.byte3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07666_ _03283_ _03285_ _03286_ _03287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_04878_ _00622_ _00031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09405_ ci_neuron.output_memory\[5\] _04628_ _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07597_ _03220_ _03221_ _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06617_ _02245_ _02202_ _02244_ _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_109_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06548_ _02086_ _02189_ _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09336_ _04099_ ci_neuron.input_memory\[1\]\[26\] _04578_ _04581_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_106_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09267_ _04537_ _04139_ _04538_ _04535_ _04539_ _00478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_23_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06479_ _00163_ _02121_ _02122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08218_ _03740_ _03742_ _03745_ _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_7_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09198_ _04499_ _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08149_ _03684_ _03686_ _03687_ _03688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_113_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10111_ _00235_ net287 ci_neuron.uut_simple_neuron.titan_id_4\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10042_ _00527_ net143 ci_neuron.output_val_internal\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08822__A2 _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09622__I1 ci_neuron.output_memory\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout290_I net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05850_ _01453_ _01489_ _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05454__I _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07520_ _03135_ _03139_ _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05781_ _01236_ _01408_ _01443_ _01444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_89_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08510__A1 ci_neuron.value_i\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07451_ _03076_ _03026_ _03077_ _03078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07382_ _03007_ _03009_ _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06402_ _01926_ _02004_ _02046_ _02047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_45_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06333_ _01943_ _01979_ _01980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_85_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09121_ ci_neuron.uut_simple_neuron.titan_id_6\[4\] _04457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_79_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06264_ _01884_ _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09052_ _04385_ _04397_ _04398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06195_ _01825_ _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05215_ _00891_ _00892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08003_ ci_neuron.uut_simple_neuron.titan_id_2\[28\] ci_neuron.uut_simple_neuron.titan_id_5\[28\]
+ _03568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05146_ _00802_ _00825_ _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09613__I1 ci_neuron.output_memory\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05077_ _00753_ _00760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09954_ _00469_ net88 ci_neuron.uut_simple_neuron.x0\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08905_ _04290_ _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09885_ _00046_ net20 ci_neuron.value_i\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08836_ _04185_ _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09392__I3 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05979_ _01593_ _01596_ _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08767_ _04216_ _00301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_28_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07718_ ci_neuron.uut_simple_neuron.titan_id_4\[13\] ci_neuron.uut_simple_neuron.titan_id_3\[13\]
+ _03330_ _03331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08698_ _04133_ _04160_ _04161_ _00287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07649_ _03225_ _03270_ _03273_ _03274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_0_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09319_ _04571_ _00498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08804__A2 _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06291__A2 _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09604__I1 ci_neuron.output_memory\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10025_ ci_neuron.input_memory\[1\]\[25\] net86 ci_neuron.uut_simple_neuron.titan_id_1\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05554__A1 _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06833__I _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05000_ _00695_ _00048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_74_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06951_ _02301_ _02307_ _02585_ _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_94_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09670_ _00257_ net260 ci_neuron.uut_simple_neuron.x3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05902_ _01538_ _01542_ _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06882_ _02515_ _02517_ _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08621_ _03879_ _04082_ _03890_ _04096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05833_ _01493_ _01494_ _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05545__A1 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Left_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05764_ _01419_ _01420_ _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08552_ _03817_ _04030_ _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07503_ _00162_ _03129_ _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08483_ ci_neuron.value_i\[5\] _03952_ _03978_ _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_07434_ _03061_ _00246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05695_ _01323_ _01348_ _01349_ _01284_ _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_85_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07365_ _02963_ _02970_ _02992_ _02993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_9_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07296_ _02862_ _02872_ _02925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06316_ _01900_ _01932_ _01962_ _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_5_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09104_ _04419_ ci_neuron.stream_o\[15\] _04445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06247_ _01880_ _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09035_ _04355_ _04382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06178_ _01826_ _01828_ _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05129_ _00773_ _00795_ _00767_ _00809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09937_ _00452_ net177 ci_neuron.uut_simple_neuron.x0\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_5_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07525__A2 _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09868_ _00059_ net29 ci_neuron.value_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08819_ _04094_ _01573_ _04246_ _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09799_ _00378_ net48 internal_ih.byte6\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09278__A2 _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07289__A1 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07461__A1 ci_neuron.uut_simple_neuron.x3\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05775__A1 _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08713__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10008_ ci_neuron.input_memory\[1\]\[8\] net204 ci_neuron.uut_simple_neuron.titan_id_1\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05480_ _01149_ _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07150_ _02780_ _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_89_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07081_ _01936_ _01868_ _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06101_ _00738_ _01751_ _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_30_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06032_ _01654_ _01678_ _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout117 net118 net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout128 net130 net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout106 net117 net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09722_ _00301_ net257 ci_neuron.uut_simple_neuron.x2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout139 net146 net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07983_ _03544_ _03548_ _03550_ _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06934_ _02526_ _02568_ _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_2_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06865_ ci_neuron.uut_simple_neuron.x3\[18\] ci_neuron.uut_simple_neuron.x3\[19\]
+ _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_87_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08555__I1 _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09653_ _04825_ _00578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05816_ ci_neuron.uut_simple_neuron.x2\[23\] _01380_ _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09584_ _04786_ _00548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08604_ _04081_ _04082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06796_ _02378_ _02397_ _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08535_ _04023_ _02226_ _03969_ _04024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05747_ _01366_ _01393_ _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05678_ _01342_ _01328_ _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08466_ _03730_ _03958_ _03953_ _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07417_ _01988_ _01958_ _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_80_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08397_ _03898_ _03901_ _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07348_ _02847_ _02975_ _02976_ _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_98_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07279_ _02897_ _02908_ _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09018_ internal_ih.data_pointer\[0\] _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07994__A2 ci_neuron.uut_simple_neuron.titan_id_5\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09196__A1 _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06182__A1 ci_neuron.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09510__I3 _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_78_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_87_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_71_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08103__I _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04980_ internal_ih.byte1\[7\] _00680_ _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06650_ _02003_ _02141_ _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_91_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05601_ _01267_ _01265_ _01268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_69_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08974__S _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06581_ _02186_ _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_87_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_96_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05532_ _01158_ _01161_ _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_82_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08320_ _03833_ _03834_ _00178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05463_ _01058_ _01132_ _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08251_ _03770_ _03772_ _03774_ _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07202_ _02789_ _02792_ _02832_ _02833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_117_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05394_ _00999_ _01066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08182_ _03715_ _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_125_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07133_ _02699_ _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07064_ _02656_ _02696_ _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07976__A2 ci_neuron.uut_simple_neuron.titan_id_5\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06015_ _01616_ _01672_ _01673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_93_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09568__I3 ci_neuron.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07966_ _03535_ _03536_ _03537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06917_ _02551_ _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08528__I1 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09705_ _00284_ net130 internal_ih.spi_rx_byte_i\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07897_ ci_neuron.uut_simple_neuron.titan_id_2\[11\] ci_neuron.uut_simple_neuron.titan_id_5\[11\]
+ _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09636_ _04810_ _04816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06848_ _02476_ _02483_ _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06779_ _02361_ _02400_ _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09567_ ci_neuron.output_memory\[29\] _04766_ _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09498_ _04697_ _04711_ _04713_ _04714_ _00534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_37_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08518_ _03945_ _04008_ _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08449_ _03941_ _03947_ _03949_ _00250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07299__I ci_neuron.uut_simple_neuron.x3\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10273_ _00566_ net153 ci_neuron.stream_o\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09019__I internal_ih.data_pointer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08858__I _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07655__A1 ci_neuron.uut_simple_neuron.titan_id_4\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07407__A1 _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout216_I net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06630__A2 _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07820_ _03415_ _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07751_ _03342_ _03343_ _03357_ _03358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06702_ _02223_ _02340_ _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_79_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04963_ _00674_ _00062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06288__I _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07682_ _03299_ _03300_ _03301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04894_ _00605_ _00633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_126_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06633_ _01994_ _02236_ _02272_ _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__08930__I1 internal_ih.byte4\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09421_ _04627_ _04643_ _04647_ _04648_ _00523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06564_ _02204_ _02205_ _02206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout31_I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09352_ _00583_ _04353_ _04589_ _00513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05515_ ci_neuron.uut_simple_neuron.x2\[17\] _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08303_ _03814_ _03819_ _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06495_ _01995_ _02097_ _02137_ _02138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09283_ _03967_ ci_neuron.input_memory\[1\]\[3\] _04543_ _04551_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05446_ _01074_ _01077_ _01115_ _01117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08234_ _03759_ _00197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_95_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05377_ _01012_ _01020_ _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08165_ ci_neuron.uut_simple_neuron.titan_id_1\[27\] ci_neuron.uut_simple_neuron.titan_id_0\[27\]
+ _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07116_ _02743_ _02747_ _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__04880__B2 _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08096_ _03644_ _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07047_ _02551_ _02624_ _02679_ _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_2_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08998_ _04348_ _00400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07949_ _03520_ _03521_ _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08921__I1 internal_ih.byte3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09619_ _04806_ _00563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07637__A1 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10256_ _00550_ net68 ci_neuron.interrupt_enabled vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10187_ _00085_ net75 ci_neuron.uut_simple_neuron.titan_id_2\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08912__I1 internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06280_ _01853_ _01906_ _01927_ _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05300_ _00973_ _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05231_ _00889_ _00899_ _00906_ _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05162_ _00813_ _00817_ _00839_ _00841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_12_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout8 net9 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_77_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05093_ _00744_ _00758_ _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09970_ _00485_ net179 ci_neuron.input_memory\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08921_ internal_ih.byte4\[5\] internal_ih.byte3\[5\] _04301_ _04305_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08852_ internal_ih.byte0\[7\] internal_ih.spi_rx_byte_i\[7\] _04264_ _04266_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07803_ _03396_ _03397_ _03400_ _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout79_I net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05995_ _01568_ _01629_ _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08783_ _04226_ _00307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07734_ _03342_ _03343_ _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04946_ _00664_ _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07665_ ci_neuron.uut_simple_neuron.titan_id_4\[4\] ci_neuron.uut_simple_neuron.titan_id_3\[4\]
+ _03286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06616_ _02241_ _02243_ _02256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04877_ internal_ih.byte7\[6\] _00616_ _00621_ _00597_ _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09404_ _04627_ _04629_ _04632_ _04634_ _00520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__05650__I _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07596_ _03152_ _03211_ _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06547_ _02186_ _02188_ _02189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_62_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09335_ _04580_ _00505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06478_ _02079_ _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09266_ spi_interface_cvonk.state\[1\] _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05429_ _00969_ _01005_ _01052_ _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_62_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08217_ _03743_ _03744_ _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09197_ _04486_ _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08148_ ci_neuron.uut_simple_neuron.titan_id_1\[24\] ci_neuron.uut_simple_neuron.titan_id_0\[24\]
+ _03687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08079_ _03627_ _03628_ _03629_ _03630_ _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_10110_ _00234_ net287 ci_neuron.uut_simple_neuron.titan_id_4\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10041_ _00526_ net143 ci_neuron.output_val_internal\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05097__A1 _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06340__B _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _00135_ net159 ci_neuron.uut_simple_neuron.titan_id_6\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout283_I net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05780_ _01411_ _01442_ _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08897__I0 internal_ih.byte3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08510__A2 _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07450_ _03004_ _03021_ _03077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06401_ _02044_ _02045_ _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07381_ _02868_ _03008_ _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08649__I0 _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06332_ _01976_ _01978_ _01979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08781__I _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09120_ _04456_ _00414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09051_ _04358_ ci_neuron.stream_o\[10\] _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_20_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06263_ _01890_ _01909_ _01911_ _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08002_ ci_neuron.uut_simple_neuron.titan_id_2\[28\] ci_neuron.uut_simple_neuron.titan_id_5\[28\]
+ _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06194_ _01820_ _01845_ _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05214_ _00811_ _00846_ ci_neuron.uut_simple_neuron.x2\[8\] _00891_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_05145_ _00782_ _00819_ _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06588__A1 _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05076_ _00737_ _00745_ _00759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09953_ _00468_ net95 ci_neuron.uut_simple_neuron.x0\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08904_ _04295_ _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09884_ _00045_ net20 ci_neuron.value_i\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08835_ _04255_ _00330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08766_ _03967_ _00758_ _04208_ _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05978_ _01634_ _01636_ _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07717_ _03326_ _03327_ _03329_ _03330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09385__S0 _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08697_ internal_ih.spi_rx_byte_i\[5\] _04148_ _04161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04929_ internal_ih.byte6\[1\] _00652_ _00653_ internal_ih.byte2\[1\] _00655_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07648_ _03271_ _03214_ _03272_ _03213_ _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_67_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07579_ _02079_ _03204_ _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_95_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09318_ _04059_ ci_neuron.input_memory\[1\]\[18\] _04567_ _04571_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06815__A2 _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09249_ _04528_ _00471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_112_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10024_ ci_neuron.input_memory\[1\]\[24\] net86 ci_neuron.uut_simple_neuron.titan_id_1\[26\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05242__A1 _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09508__A1 ci_neuron.output_memory\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06950_ _02578_ _02584_ _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06881_ _02422_ _02460_ _02516_ _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05901_ _01523_ _01537_ _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input3_I spi_pico_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05832_ _01448_ _01451_ _01491_ _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08620_ _04095_ _00275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05763_ _01421_ _01424_ _01386_ _01425_ _01343_ _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_08551_ _03809_ _04036_ _03825_ _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05694_ _01358_ _00212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07502_ _03126_ _03128_ _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08482_ _03965_ _03976_ _03977_ _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_07433_ _02990_ _03060_ _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_85_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07364_ _02966_ _02969_ _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout8_I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09103_ _04415_ _04443_ _04444_ _00409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07295_ _02879_ _02883_ _02923_ _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06315_ _01959_ _01961_ _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06246_ _01894_ _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_103_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09034_ _04370_ _04381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_107_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06177_ _01829_ _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05128_ _00787_ _00807_ _00808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05059_ _00743_ _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09936_ _00451_ net177 ci_neuron.uut_simple_neuron.x0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09867_ _00058_ net28 ci_neuron.value_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06733__A1 _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07590__I _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_116_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08818_ _04224_ _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09798_ _00377_ net41 internal_ih.byte5\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08749_ _04194_ _04203_ _00296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08635__B _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09310__I _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_125_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07461__A2 ci_neuron.uut_simple_neuron.x3\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10007_ ci_neuron.input_memory\[1\]\[7\] net204 ci_neuron.uut_simple_neuron.titan_id_1\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_125_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08477__A1 _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07080_ _02710_ _02711_ _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06100_ _01755_ _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06031_ _01648_ _01681_ _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05463__A1 _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout118 net119 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout107 net111 net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout129 net130 net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07982_ _03545_ _03550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06933_ _02528_ _02567_ _02568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06963__A1 _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09721_ _00300_ net256 ci_neuron.uut_simple_neuron.x2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_2_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06864_ _02383_ _02448_ _02499_ _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout61_I net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09652_ ci_neuron.stream_o\[27\] ci_neuron.output_memory\[27\] _04821_ _04825_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06795_ _02378_ _02397_ _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05815_ _01474_ _01476_ _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09583_ _04605_ ci_neuron.normalised_stream_write_address\[0\] _04785_ _04786_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08603_ _03863_ _04077_ _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05746_ _01366_ _01393_ _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08534_ _04020_ _04022_ _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_38_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08468__A1 ci_neuron.value_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05677_ ci_neuron.uut_simple_neuron.x2\[21\] _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08465_ _03729_ _03958_ _03963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07416_ _03042_ _03043_ _03044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08396_ _03895_ _03899_ _03900_ _03894_ _03901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07347_ _02850_ _02909_ _02976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_98_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07278_ _02899_ _02907_ _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09017_ _04355_ _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06229_ _01873_ _01878_ _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09919_ _00016_ net8 ci_neuron.address_i\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08631__A1 _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07198__A1 _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05600_ _01226_ _01264_ _01267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_69_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06580_ _02191_ _02194_ _02220_ _02221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_91_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05531_ _01166_ _01199_ _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_82_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05462_ _01106_ _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08250_ _03773_ _03766_ _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07201_ _02821_ _02831_ _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_15_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08181_ _03707_ _03713_ _03712_ _03703_ _03714_ _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_07132_ _02761_ _02763_ _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_05393_ _00932_ _01064_ _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07063_ _02658_ _02695_ _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_113_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06014_ _01666_ _01671_ _01672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07965_ ci_neuron.uut_simple_neuron.titan_id_2\[23\] ci_neuron.uut_simple_neuron.titan_id_5\[23\]
+ _03536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06916_ ci_neuron.uut_simple_neuron.x3\[19\] _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09704_ _00283_ net128 internal_ih.spi_rx_byte_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09635_ _04815_ _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07896_ _03478_ _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06847_ _02479_ _02482_ _02483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06778_ _02415_ _00236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09566_ _04765_ _04767_ _04770_ _04772_ _00544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05729_ _01388_ _01392_ _01393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09497_ ci_neuron.output_val_internal\[18\] _04705_ _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08517_ _04006_ _04007_ _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08448_ _02898_ _03948_ _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08379_ _03882_ _03876_ _03885_ _03881_ _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_60_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10272_ _00565_ net154 ci_neuron.stream_o\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09495__I3 _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout111_I net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08114__I _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout209_I net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06394__A2 _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07750_ ci_neuron.uut_simple_neuron.titan_id_4\[16\] ci_neuron.uut_simple_neuron.titan_id_3\[16\]
+ _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04962_ internal_ih.byte0\[7\] _00670_ _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06701_ _02337_ _02339_ _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_07681_ ci_neuron.uut_simple_neuron.titan_id_4\[7\] ci_neuron.uut_simple_neuron.titan_id_3\[7\]
+ _03300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04893_ _00632_ _00018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06632_ _01995_ _02135_ _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09420_ ci_neuron.output_val_internal\[7\] _04633_ _04648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06563_ _02160_ _02158_ _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09351_ _04145_ _04152_ _04352_ _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_47_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05514_ _01175_ _01182_ _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09282_ _03961_ _04544_ _04550_ _00482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08302_ _03816_ _03818_ _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_118_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06494_ _02135_ _02136_ _02137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_75_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08233_ _03754_ _03756_ _03758_ _03759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05445_ _01074_ _01077_ _01115_ _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_43_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05376_ _00860_ _01044_ _01047_ _01048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_7_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08164_ _03693_ _03698_ _03700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07115_ _02225_ _02746_ _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_95_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08095_ ci_neuron.uut_simple_neuron.titan_id_1\[15\] ci_neuron.uut_simple_neuron.titan_id_0\[15\]
+ _03644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07046_ _02555_ _02623_ _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08997_ internal_ih.current_instruction\[6\] _04341_ _04348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_98_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07948_ _03517_ _03518_ _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07879_ ci_neuron.uut_simple_neuron.titan_id_2\[8\] ci_neuron.uut_simple_neuron.titan_id_5\[8\]
+ _03461_ _03462_ _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09618_ ci_neuron.stream_o\[12\] ci_neuron.output_memory\[12\] _04805_ _04806_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_104_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09549_ ci_neuron.output_val_internal\[26\] _04749_ _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09011__A1 internal_ih.data_pointer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10255_ _00549_ net105 ci_neuron.normalised_stream_write_address\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10186_ _00084_ net75 ci_neuron.uut_simple_neuron.titan_id_2\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout290 net291 net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07325__A1 _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__A2 ci_neuron.uut_simple_neuron.titan_id_5\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07013__I _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08109__I _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05230_ _00890_ _00898_ _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_25_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05161_ _00813_ _00817_ _00839_ _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_71_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout9 net18 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05092_ _00773_ _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08920_ _04304_ _00366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10026__D ci_neuron.input_memory\[1\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08851_ _04265_ _00336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07802_ ci_neuron.uut_simple_neuron.titan_id_4\[27\] ci_neuron.uut_simple_neuron.titan_id_3\[27\]
+ _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05994_ _01649_ _01651_ _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08782_ _04003_ _00896_ _04225_ _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07733_ ci_neuron.uut_simple_neuron.titan_id_4\[16\] ci_neuron.uut_simple_neuron.titan_id_3\[16\]
+ _03343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04945_ _00599_ _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07664_ ci_neuron.uut_simple_neuron.titan_id_4\[4\] ci_neuron.uut_simple_neuron.titan_id_3\[4\]
+ _03285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07867__A2 ci_neuron.uut_simple_neuron.titan_id_5\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04876_ internal_ih.byte4\[6\] internal_ih.byte3\[6\] _00601_ _00621_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06615_ _02247_ _02255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09403_ ci_neuron.output_val_internal\[4\] _04633_ _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07595_ _03155_ _03210_ _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06546_ _02094_ _02187_ _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08816__A1 _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09334_ _04094_ ci_neuron.input_memory\[1\]\[25\] _04578_ _04580_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06477_ _02113_ _02063_ _02112_ _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09265_ _04166_ _04138_ _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05428_ _00939_ _01054_ _01091_ _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_63_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09196_ _03974_ _04494_ _04498_ _00448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08216_ _03733_ _03737_ _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05359_ _01004_ _01022_ _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_15_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08147_ ci_neuron.uut_simple_neuron.titan_id_1\[24\] ci_neuron.uut_simple_neuron.titan_id_0\[24\]
+ _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08078_ ci_neuron.uut_simple_neuron.titan_id_1\[11\] ci_neuron.uut_simple_neuron.titan_id_0\[11\]
+ _03630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07029_ _02178_ _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_101_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10040_ _00525_ net143 ci_neuron.output_val_internal\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07307__A1 _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09480__A1 ci_neuron.output_memory\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05097__A2 _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10238_ _00134_ net191 ci_neuron.uut_simple_neuron.titan_id_6\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10169_ _00095_ net210 ci_neuron.uut_simple_neuron.titan_id_2\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_128_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout276_I net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09223__I _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06400_ _02003_ _02045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07380_ ci_neuron.uut_simple_neuron.x3\[26\] ci_neuron.uut_simple_neuron.x3\[27\]
+ _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08649__I1 ci_neuron.uut_simple_neuron.x3\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06331_ _01890_ _01944_ _01917_ _01977_ _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_84_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06262_ _01827_ _01884_ _01910_ _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_79_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09050_ _04378_ _04395_ _04396_ _00404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05213_ _00742_ _00862_ _00870_ _00890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08001_ _03566_ _00147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06193_ _01842_ _01844_ _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_111_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05144_ _00810_ _00823_ _00824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06588__A2 _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05075_ _00757_ _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout91_I net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09952_ _00467_ net95 ci_neuron.uut_simple_neuron.x0\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08903_ internal_ih.byte3\[5\] internal_ih.byte2\[5\] _04291_ _04295_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09883_ _00043_ net23 ci_neuron.value_i\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08834_ internal_ih.byte0\[0\] _04143_ _04254_ _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08765_ _03961_ _04209_ _04215_ _00300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05977_ _01076_ _01592_ _01635_ _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07716_ ci_neuron.uut_simple_neuron.titan_id_4\[12\] ci_neuron.uut_simple_neuron.titan_id_3\[12\]
+ _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_68_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09385__S1 _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08696_ internal_ih.spi_tx_byte_o\[4\] _04136_ _04157_ internal_ih.spi_rx_byte_i\[4\]
+ _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_04928_ _00654_ _00008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07647_ _03146_ _03143_ _03272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04859_ internal_ih.byte4\[1\] internal_ih.byte3\[1\] _00608_ _00609_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_0_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07578_ _02088_ _02103_ _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06529_ _02130_ _02151_ _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09317_ _04570_ _00497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09248_ _04104_ _03892_ _04525_ _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_105_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09179_ _04485_ _04206_ _04486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09517__A2 _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10023_ ci_neuron.input_memory\[1\]\[23\] net95 ci_neuron.uut_simple_neuron.titan_id_1\[25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09043__I internal_ih.data_pointer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09453__A1 ci_neuron.output_memory\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09205__A1 _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06880_ _02424_ _02459_ _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05900_ _01389_ _01558_ _01559_ _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05831_ _01492_ _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05762_ _00749_ _01384_ _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08550_ _04030_ _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07501_ _02074_ _03127_ _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05693_ _01355_ _01357_ _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08481_ _03739_ _03963_ _03741_ _03977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07432_ _02991_ _03059_ _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_85_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08792__I _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07363_ _02974_ _02977_ _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09102_ internal_ih.spi_tx_byte_o\[6\] _04427_ _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_128_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07294_ _02856_ _02853_ _02878_ _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06314_ _01960_ _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06245_ _01891_ _01893_ _01894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09033_ _04372_ _04378_ _04380_ _00403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06176_ _01819_ _01828_ _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07758__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05127_ _00792_ _00797_ _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05058_ _00742_ _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09935_ _00450_ net177 ci_neuron.uut_simple_neuron.x0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09866_ _00055_ net28 ci_neuron.value_i\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08817_ _01473_ _04236_ _04245_ _00322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08183__A1 _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09797_ _00376_ net41 internal_ih.byte5\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08748_ internal_ih.received_byte_count\[6\] _04202_ _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_95_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08486__A2 _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08679_ spi_interface_cvonk.SS_r\[1\] _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_83_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08797__I0 _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08877__I _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10006_ ci_neuron.input_memory\[1\]\[6\] net206 ci_neuron.uut_simple_neuron.titan_id_1\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_125_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06724__A2 _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09501__I _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06030_ _01652_ _01680_ _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08788__I0 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout119 net217 net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout108 net111 net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07981_ _03549_ _00144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06932_ _02538_ _02540_ _02566_ _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09720_ _00299_ net219 ci_neuron.uut_simple_neuron.x2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_2_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04974__A1 internal_ih.byte1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06863_ _02388_ _02498_ _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_87_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09651_ _04824_ _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06794_ _02365_ _02430_ _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05814_ _00748_ _01475_ _01476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08602_ _03986_ _04079_ _04080_ _00272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09582_ _04599_ _00730_ _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05745_ _01406_ _01407_ _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08533_ _03789_ _04006_ _04021_ _03959_ _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_38_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06479__A1 _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08468__A2 _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05676_ _01338_ _01340_ _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08464_ _03957_ _03961_ _03962_ _00252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07415_ _02953_ _02959_ _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08395_ ci_neuron.uut_simple_neuron.x0\[26\] _03891_ _03900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07346_ _02850_ _02909_ _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07277_ _02902_ _02906_ _02907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_60_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09016_ _04358_ ci_neuron.stream_o\[0\] ci_neuron.stream_o\[16\] _04359_ _04363_
+ _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_33_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06228_ ci_neuron.uut_simple_neuron.x3\[5\] _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06159_ ci_neuron.uut_simple_neuron.x2\[31\] _01812_ _01813_ _01814_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09918_ _00015_ net6 ci_neuron.address_i\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04965__A1 internal_ih.byte1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08156__A1 _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09849_ _00428_ net158 ci_neuron.output_memory\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08631__A2 _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04956__A1 internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05920__A3 _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05530_ _01124_ _01198_ _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_82_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05461_ _01088_ _01095_ _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07200_ _02824_ _02830_ _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05392_ _01032_ _01063_ _01064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08180_ ci_neuron.uut_simple_neuron.titan_id_1\[29\] ci_neuron.uut_simple_neuron.titan_id_0\[29\]
+ _03714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07131_ _02649_ _02698_ _02762_ _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10029__D ci_neuron.input_memory\[1\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08083__B1 _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07062_ _02668_ _02694_ _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06013_ _00936_ _01668_ _01670_ _01671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05934__I _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04947__A1 internal_ih.byte0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07964_ _03533_ _03534_ _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06915_ _02380_ _02503_ _02549_ _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07895_ ci_neuron.uut_simple_neuron.titan_id_2\[11\] ci_neuron.uut_simple_neuron.titan_id_5\[11\]
+ _03477_ _03478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09703_ _00282_ net121 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06846_ _01824_ _02481_ _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09634_ ci_neuron.stream_o\[19\] ci_neuron.output_memory\[19\] _04811_ _04815_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06777_ _02410_ _02414_ _02415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05372__A1 _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09565_ ci_neuron.output_val_internal\[28\] _04771_ _04772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08466__B _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05728_ _01389_ _01391_ _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08516_ _03782_ _03997_ _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09496_ _04701_ _04712_ _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05659_ _01146_ _01223_ _01287_ _01324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_08447_ _03940_ _03948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08378_ _03874_ _03875_ _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07329_ _01968_ _02957_ _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10271_ _00564_ net154 ci_neuron.stream_o\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08924__I0 internal_ih.byte4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09252__S _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05363__A1 _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout90 net91 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09652__I1 ci_neuron.output_memory\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05418__A2 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout104_I net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06918__A2 _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04929__B2 internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04961_ _00673_ _00061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06700_ _02283_ _02338_ _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07680_ _03295_ _03297_ _03298_ _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_04892_ internal_ih.byte4\[3\] _00625_ _00628_ internal_ih.byte0\[3\] _00632_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06631_ _02219_ _02269_ _02270_ _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06562_ _02154_ _02157_ _02204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09350_ _04588_ _00512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05513_ _01179_ _01181_ _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09281_ ci_neuron.input_memory\[1\]\[2\] _04549_ _04550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08301_ _03811_ _03817_ _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_19_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06493_ _02096_ _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08232_ _03742_ _03754_ _03757_ _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05444_ _01078_ _01114_ _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout17_I net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05375_ _01017_ _01046_ _01047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09643__I1 ci_neuron.output_memory\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08163_ _03699_ _00083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07114_ _02234_ _02745_ _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_95_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08094_ _03639_ _03640_ _03642_ _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_31_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07045_ _02495_ _02626_ _02677_ _02678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_42_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_10_Left_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08996_ _04347_ _00399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07582__A2 _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07947_ ci_neuron.uut_simple_neuron.titan_id_2\[20\] ci_neuron.uut_simple_neuron.titan_id_5\[20\]
+ _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08531__A1 ci_neuron.value_i\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07878_ _03463_ _00157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06829_ _02463_ _02465_ _02466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09617_ _04789_ _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_104_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09548_ _04746_ _04756_ _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09479_ _04674_ _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06845__A1 _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04856__B1 _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09634__I1 ci_neuron.output_memory\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09011__A2 internal_ih.data_pointer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10254_ _00548_ net105 ci_neuron.normalised_stream_write_address\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10185_ _00083_ net80 ci_neuron.uut_simple_neuron.titan_id_2\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout291 net4 net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout280 net281 net280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08522__A1 _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05336__A1 _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05749__I _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05160_ _00733_ _00835_ _00838_ _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08589__A1 _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05091_ _00760_ _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09002__A2 _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08850_ internal_ih.byte0\[6\] internal_ih.spi_rx_byte_i\[6\] _04264_ _04265_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07801_ ci_neuron.uut_simple_neuron.titan_id_4\[28\] ci_neuron.uut_simple_neuron.titan_id_3\[28\]
+ _03399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07564__A2 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08761__A1 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05993_ _01650_ _01631_ _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08781_ _04224_ _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07732_ _03338_ _03340_ _03341_ _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_04944_ _00663_ _00016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05327__A1 _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07663_ _03284_ _00120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04875_ _00620_ _00030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06614_ _02254_ _00233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09402_ _04610_ _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07594_ _02808_ _03217_ _03218_ _03219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_75_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09333_ _04579_ _00504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06545_ ci_neuron.uut_simple_neuron.x3\[12\] ci_neuron.uut_simple_neuron.x3\[13\]
+ _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08816__A2 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06476_ _02070_ _02116_ _02118_ _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09264_ spi_interface_cvonk.state\[1\] _04127_ _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05427_ _01097_ _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08215_ _03730_ _03740_ _03743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09195_ _03740_ _04491_ _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08146_ _03685_ _00080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05358_ _01004_ _01022_ _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07252__A1 _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05289_ ci_neuron.uut_simple_neuron.x2\[9\] _00910_ ci_neuron.uut_simple_neuron.x2\[11\]
+ _00963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08077_ ci_neuron.uut_simple_neuron.titan_id_1\[11\] ci_neuron.uut_simple_neuron.titan_id_0\[11\]
+ ci_neuron.uut_simple_neuron.titan_id_1\[10\] ci_neuron.uut_simple_neuron.titan_id_0\[10\]
+ _03629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_07028_ _01846_ _02659_ _02660_ _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08979_ _04337_ _00392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09741__D _00320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09304__I0 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06953__I _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_117_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10237_ _00133_ net208 ci_neuron.uut_simple_neuron.titan_id_6\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10168_ _00094_ net210 ci_neuron.uut_simple_neuron.titan_id_2\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_128_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10099_ _00165_ net274 ci_neuron.uut_simple_neuron.titan_id_4\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout171_I net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06330_ _01940_ _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06261_ _01871_ _01883_ _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_79_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05212_ _00835_ _00888_ _00869_ _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08000_ ci_neuron.uut_simple_neuron.titan_id_2\[28\] ci_neuron.uut_simple_neuron.titan_id_5\[28\]
+ _03565_ _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06192_ ci_neuron.uut_simple_neuron.x3\[1\] _01843_ _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_13_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05143_ _00818_ _00819_ _00822_ _00784_ _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05074_ _00756_ _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09951_ _00466_ net82 ci_neuron.uut_simple_neuron.x0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08982__A1 _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08902_ _04294_ _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09882_ _00042_ net23 ci_neuron.value_i\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05548__A1 _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08833_ _04192_ _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05976_ _01556_ _01591_ _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08764_ _00774_ _04214_ _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07715_ _03328_ _00098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04927_ internal_ih.byte6\[0\] _00652_ _00653_ internal_ih.byte2\[0\] _00654_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08695_ _04134_ _04158_ _04159_ _00286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07646_ _03066_ _03141_ _03271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_94_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04858_ _00600_ _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_0_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07577_ _03201_ _03202_ _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06528_ _02168_ _02169_ _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09316_ _04052_ ci_neuron.input_memory\[1\]\[17\] _04567_ _04570_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09247_ _04527_ _00470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09462__A2 _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06459_ _02102_ _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09178_ _03934_ _03936_ _04485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08129_ _03668_ _03669_ _03671_ _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_31_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10022_ ci_neuron.input_memory\[1\]\[22\] net93 ci_neuron.uut_simple_neuron.titan_id_1\[24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05830_ _01448_ _01451_ _01491_ _01492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07500_ _02081_ _02480_ _03127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05761_ _01105_ _01422_ _01371_ _01373_ _01423_ _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05692_ _01304_ _01314_ _01356_ _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08480_ _03739_ _03741_ _03963_ _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_07431_ _02993_ _03055_ _03058_ _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_92_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07362_ _02988_ _02989_ _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06313_ ci_neuron.uut_simple_neuron.x3\[7\] _01960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09101_ ci_neuron.stream_o\[30\] _04416_ _04442_ _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07293_ _02885_ _02895_ _02921_ _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06244_ _01892_ _01841_ _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09032_ internal_ih.spi_tx_byte_o\[0\] _04379_ _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06175_ ci_neuron.uut_simple_neuron.x3\[1\] ci_neuron.uut_simple_neuron.x3\[2\] _01828_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05126_ _00804_ _00805_ _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_111_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05057_ _00741_ _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09934_ _00449_ net177 ci_neuron.uut_simple_neuron.x0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_09865_ _00044_ net28 ci_neuron.value_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08816_ _04089_ _04237_ _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_5_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07930__A2 ci_neuron.uut_simple_neuron.titan_id_5\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09796_ _00375_ net39 internal_ih.byte5\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05959_ _01472_ _01532_ _01579_ _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08747_ _04193_ _04201_ _04202_ _00295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_95_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08678_ _04145_ _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07629_ _03252_ _03253_ _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06497__A2 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_2_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_39_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10005_ ci_neuron.input_memory\[1\]\[5\] net202 ci_neuron.uut_simple_neuron.titan_id_1\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_125_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07988__A2 ci_neuron.uut_simple_neuron.titan_id_5\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_57_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout109 net111 net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07980_ _03546_ _03548_ _03549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06931_ _02544_ _02565_ _02566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09650_ ci_neuron.stream_o\[26\] ci_neuron.output_memory\[26\] _04821_ _04824_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06862_ ci_neuron.uut_simple_neuron.x3\[18\] _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_87_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08601_ _02805_ _04011_ _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06793_ _02427_ _02429_ _02430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05813_ ci_neuron.uut_simple_neuron.x2\[24\] _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_66_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09581_ _04765_ _04781_ _04783_ _04784_ _00547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05744_ _00934_ _01395_ _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08532_ _03799_ _04006_ _04021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06479__A2 _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08463_ _01849_ _03948_ _03962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07414_ _02956_ _02958_ _03042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05675_ _01186_ _01287_ _01339_ _01146_ _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_65_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07212__I _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08394_ _03889_ _03891_ _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_128_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07345_ _02973_ _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07276_ _02904_ _02905_ _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06227_ _01876_ _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09015_ _04360_ _04362_ _04363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06158_ _01464_ _01462_ _01454_ _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06089_ _01700_ _01719_ _01745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05109_ _00780_ _00782_ _00783_ _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_111_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09917_ _00014_ net8 ci_neuron.address_i\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09848_ _00427_ net191 ci_neuron.output_memory\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05914__A1 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09779_ _00358_ net63 internal_ih.byte3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout251_I net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05460_ _01129_ _01095_ _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05391_ _01034_ _01038_ _01062_ _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_15_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07130_ _02652_ _02697_ _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07061_ _02671_ _02693_ _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_100_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06012_ _00738_ _01669_ _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07963_ _03530_ _03531_ _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06914_ _02547_ _02548_ _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06149__A1 _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_74_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07894_ _03473_ _03474_ _03476_ _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09702_ spi_interface_cvonk.MOSI_r\[0\] net128 internal_ih.spi_rx_byte_i\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06845_ _02038_ _02480_ _02481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09633_ _04814_ _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09564_ _04704_ _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06776_ _02308_ _02412_ _02413_ _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08515_ _04005_ _03998_ _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05727_ _00864_ _01207_ _01390_ _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_65_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09495_ _03841_ ci_neuron.input_memory\[1\]\[18\] _01227_ _02616_ _04691_ _04692_
+ _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_05658_ _01321_ _01295_ _01322_ _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_65_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08446_ ci_neuron.value_i\[0\] _03944_ _03946_ _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_93_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_83_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08377_ _03884_ _00185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07328_ _02374_ _02395_ _02957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05589_ _01255_ _01220_ _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_61_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07259_ _02282_ _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07821__A1 ci_neuron.uut_simple_neuron.titan_id_4\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10270_ _00563_ net153 ci_neuron.stream_o\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_92_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout91 net96 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_12_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04874__B2 _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout80 net83 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08860__I0 internal_ih.byte1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08612__S _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05100__I net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09565__A1 ci_neuron.output_val_internal\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04960_ internal_ih.byte0\[6\] _00670_ _00673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08915__I1 internal_ih.byte3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06630_ _02221_ _02239_ _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04891_ _00631_ _00017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06561_ _02199_ _02202_ _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06303__A1 _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06492_ _02093_ _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05512_ _01147_ _01180_ _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09280_ _04545_ _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08300_ _03808_ _03810_ _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05443_ _01081_ _01113_ _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08231_ _03748_ _03749_ _03747_ _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06854__A2 _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05374_ _00982_ _01045_ _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_70_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08162_ _03697_ _03698_ _03699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07113_ _02379_ _02685_ _02744_ _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_95_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08093_ ci_neuron.uut_simple_neuron.titan_id_1\[14\] ci_neuron.uut_simple_neuron.titan_id_0\[14\]
+ _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07044_ _02622_ _02676_ _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_70_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09417__I _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07031__A2 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08995_ internal_ih.current_instruction\[5\] _04340_ _04347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07946_ _03519_ _00139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07877_ _03461_ _03462_ _03463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08531__A2 _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06828_ _02408_ _02405_ _02464_ _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_97_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09616_ _04804_ _00562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06759_ _02393_ _02396_ _02397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_104_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09547_ _03890_ ci_neuron.input_memory\[1\]\[26\] _01579_ _03083_ _04738_ _04739_
+ _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_93_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09478_ _04696_ _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04856__A1 _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08429_ ci_neuron.address_i\[0\] _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10253_ _00151_ net44 ci_neuron.uut_simple_neuron.titan_id_6\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10184_ _00082_ net80 ci_neuron.uut_simple_neuron.titan_id_2\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout281 net282 net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout270 net271 net270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08522__A2 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08286__A1 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08589__A2 _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout214_I net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05090_ _00763_ _00771_ _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_122_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04870__I1 internal_ih.byte3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07800_ _03398_ _00114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08780_ _04207_ _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_127_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07731_ ci_neuron.uut_simple_neuron.titan_id_4\[15\] ci_neuron.uut_simple_neuron.titan_id_3\[15\]
+ _03341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05992_ _01604_ _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04943_ internal_ih.byte6\[7\] _00658_ _00659_ internal_ih.byte2\[7\] _00663_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07662_ ci_neuron.uut_simple_neuron.titan_id_4\[4\] ci_neuron.uut_simple_neuron.titan_id_3\[4\]
+ _03283_ _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_04874_ internal_ih.byte7\[5\] _00616_ _00619_ _00597_ _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06613_ _02250_ _02253_ _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07593_ _02933_ _03012_ _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09401_ _04630_ _04631_ _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06544_ _02091_ _02143_ _02185_ _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09332_ _04089_ ci_neuron.input_memory\[1\]\[24\] _04578_ _04579_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06475_ _02072_ _02115_ _02118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_75_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09263_ _04127_ _04535_ _04536_ _00477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05426_ _01096_ _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08214_ _03741_ _03742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09194_ _03734_ _04489_ _04497_ _00447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05357_ _00996_ _01025_ _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08145_ ci_neuron.uut_simple_neuron.titan_id_1\[24\] ci_neuron.uut_simple_neuron.titan_id_0\[24\]
+ _03684_ _03685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_15_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05288_ _00961_ _00892_ _00942_ _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__05263__A1 _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08076_ _03619_ _03624_ _03628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07027_ _02128_ _02603_ _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08978_ internal_ih.byte7\[6\] internal_ih.byte6\[6\] _04257_ _04337_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07929_ _03498_ _03503_ _03505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_97_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06190__B _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05585__I _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10236_ _00132_ net212 ci_neuron.uut_simple_neuron.titan_id_6\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10143__D _00208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05006__A1 internal_ih.byte3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10167_ _00093_ net210 ci_neuron.uut_simple_neuron.titan_id_2\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08896__I _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10098_ _00164_ net273 ci_neuron.uut_simple_neuron.titan_id_4\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout164_I net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06809__A2 _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06260_ _01895_ _01899_ _01908_ _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_115_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05211_ _00887_ _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_79_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06191_ ci_neuron.uut_simple_neuron.x3\[2\] _01838_ _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08806__I0 _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08580__B _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05142_ _00821_ _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05073_ ci_neuron.uut_simple_neuron.x2\[3\] _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09950_ _00465_ net107 ci_neuron.uut_simple_neuron.x0\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08982__A2 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08901_ internal_ih.byte3\[4\] internal_ih.byte2\[4\] _04291_ _04294_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_110_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09881_ _00041_ net24 ci_neuron.value_i\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08832_ _04253_ _00329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05975_ _01449_ _01633_ _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08763_ _04210_ _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07714_ _03326_ _03327_ _03328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08498__A1 _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04926_ _00626_ _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08694_ internal_ih.spi_rx_byte_i\[4\] _04149_ _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07645_ _03239_ _03260_ _03269_ _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_95_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04857_ _00607_ _00025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07576_ _02074_ _03127_ _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06527_ _01831_ _02129_ _02169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09315_ _04569_ _00496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06458_ _02100_ _02101_ _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09246_ _04099_ _03890_ _04525_ _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05409_ _01038_ _01062_ _01080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06389_ _01993_ _02011_ _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09177_ _00587_ _04187_ _04189_ _04353_ _00443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08128_ ci_neuron.uut_simple_neuron.titan_id_1\[20\] ci_neuron.uut_simple_neuron.titan_id_0\[20\]
+ _03671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08059_ _03613_ _00093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10021_ ci_neuron.input_memory\[1\]\[21\] net93 ci_neuron.uut_simple_neuron.titan_id_1\[23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09340__I _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05475__A1 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10219_ _00116_ net75 ci_neuron.uut_simple_neuron.titan_id_5\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05760_ _01375_ _01337_ _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05691_ _01300_ _01303_ _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07430_ _02918_ _03056_ _03057_ _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_85_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07361_ _02979_ _02984_ _02989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06312_ _01903_ _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09100_ _04356_ _04439_ _04441_ _04411_ _04442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07292_ _02855_ _02884_ _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09031_ _04377_ _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06243_ _01820_ _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06174_ _01826_ _01827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_53_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05125_ _00778_ _00800_ _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05056_ _00740_ _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09933_ _00448_ net171 ci_neuron.uut_simple_neuron.x0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_09864_ _00033_ net28 ci_neuron.value_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08815_ _04244_ _00321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_5_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09425__I _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09795_ _00374_ net55 internal_ih.byte5\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05958_ ci_neuron.uut_simple_neuron.x2\[1\] _01581_ _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08746_ internal_ih.received_byte_count\[5\] internal_ih.received_byte_count\[4\]
+ _04199_ _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_95_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05889_ _01547_ _01549_ _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08677_ internal_ih.spi_rx_byte_i\[1\] _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04909_ internal_ih.byte5\[1\] _00640_ _00641_ internal_ih.byte1\[1\] _00643_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07628_ _03194_ _03209_ _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07559_ _02504_ _03101_ _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09229_ _04517_ _00462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10004_ ci_neuron.input_memory\[1\]\[4\] net201 ci_neuron.uut_simple_neuron.titan_id_1\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_125_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_103_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05696__A1 _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_112_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06930_ _02546_ _02564_ _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input1_I spi_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06861_ _02330_ _02450_ _02496_ _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_87_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08600_ ci_neuron.value_i\[22\] _03971_ _04078_ _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XPHY_EDGE_ROW_121_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06792_ _01892_ _02428_ _02429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05812_ _00739_ _01473_ _01474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09580_ ci_neuron.output_val_internal\[31\] _04771_ _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05743_ _01359_ _01394_ _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08531_ ci_neuron.value_i\[12\] _04019_ _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05674_ _01223_ _01267_ _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08462_ ci_neuron.value_i\[2\] _03944_ _03960_ _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07413_ _02967_ _02968_ _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05687__A1 _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08393_ ci_neuron.uut_simple_neuron.x0\[27\] ci_neuron.uut_simple_neuron.x0\[28\]
+ _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07344_ _02918_ _02920_ _02972_ _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_18_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07275_ _01929_ _01937_ _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_98_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06226_ _01849_ _01859_ _01875_ _01876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04852__I _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09014_ _04361_ ci_neuron.stream_o\[8\] _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06157_ _01810_ _01811_ _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06088_ _01705_ _01718_ _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05108_ _00787_ _00770_ _00788_ _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09916_ _00013_ net6 ci_neuron.address_i\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05039_ _00724_ _00725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09847_ _00426_ net196 ci_neuron.output_memory\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05914__A2 _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09778_ _00357_ net63 internal_ih.byte3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08729_ _04187_ _04188_ _00587_ _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_107_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05602__A1 _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07355__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05390_ _01048_ _01051_ _01061_ _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_6_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08607__A1 _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07060_ _02688_ _02692_ _02693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06011_ ci_neuron.uut_simple_neuron.x2\[27\] ci_neuron.uut_simple_neuron.x2\[28\]
+ _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05841__A1 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06397__A2 _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09701_ net3 net128 spi_interface_cvonk.MOSI_r\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07962_ ci_neuron.uut_simple_neuron.titan_id_2\[22\] ci_neuron.uut_simple_neuron.titan_id_5\[22\]
+ _03533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06913_ _02502_ _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07893_ ci_neuron.uut_simple_neuron.titan_id_2\[10\] ci_neuron.uut_simple_neuron.titan_id_5\[10\]
+ _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06844_ _02057_ _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09632_ ci_neuron.stream_o\[18\] ci_neuron.output_memory\[18\] _04811_ _04814_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09563_ _04768_ _04769_ _04770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06775_ _02411_ _02356_ _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08514_ ci_neuron.uut_simple_neuron.x0\[10\] _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05726_ _01338_ _01340_ _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09494_ ci_neuron.output_memory\[18\] _04698_ _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05657_ _01288_ _01294_ _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_65_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08445_ _03725_ _03945_ _03946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05588_ _01254_ _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08376_ _03880_ _03883_ _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07327_ _02954_ _02955_ _02956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04883__A2 _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07258_ _02886_ _02887_ _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07189_ _02815_ _02819_ _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06209_ ci_neuron.uut_simple_neuron.x3\[2\] _01859_ _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_14_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09574__A2 _04778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout92 net94 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout70 net71 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout81 net83 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05588__I _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08860__I1 internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07308__I ci_neuron.uut_simple_neuron.x3\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07328__A1 _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04890_ internal_ih.byte4\[2\] _00625_ _00628_ internal_ih.byte0\[2\] _00631_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_126_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07879__A2 ci_neuron.uut_simple_neuron.titan_id_5\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06560_ _02200_ _02201_ _02202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_48_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06491_ _02099_ _02104_ _02133_ _02134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05511_ _01098_ _01150_ _01180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05442_ _01082_ _01112_ _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08230_ _03755_ _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05373_ _00939_ _01007_ _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08161_ ci_neuron.uut_simple_neuron.titan_id_1\[27\] ci_neuron.uut_simple_neuron.titan_id_0\[27\]
+ _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07112_ _02380_ _02547_ _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_95_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08092_ _03641_ _00069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07043_ _02552_ _02624_ _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08994_ _04346_ _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07319__A1 _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07945_ _03517_ _03518_ _03519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07876_ ci_neuron.uut_simple_neuron.titan_id_2\[8\] ci_neuron.uut_simple_neuron.titan_id_5\[8\]
+ _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09615_ ci_neuron.stream_o\[11\] ci_neuron.output_memory\[11\] _04800_ _04804_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06827_ _02401_ _02404_ _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06758_ _02395_ _02396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_92_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09546_ ci_neuron.output_memory\[26\] _04744_ _04755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05709_ _01145_ _01333_ _01372_ _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_66_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09477_ _04596_ _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06689_ _02289_ _02292_ _02327_ _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_66_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08428_ _00724_ _03924_ _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08359_ _03868_ _00183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05805__A1 _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10252_ _00150_ net45 ci_neuron.uut_simple_neuron.titan_id_6\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10183_ _00081_ net83 ci_neuron.uut_simple_neuron.titan_id_2\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout282 net283 net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout260 net262 net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout271 net272 net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_17_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06297__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07730_ ci_neuron.uut_simple_neuron.titan_id_4\[15\] ci_neuron.uut_simple_neuron.titan_id_3\[15\]
+ _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05991_ _01607_ _01630_ _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04942_ _00662_ _00015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07661_ _03279_ _03281_ _03282_ _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_04873_ internal_ih.byte4\[5\] internal_ih.byte3\[5\] _00601_ _00619_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06612_ _02166_ _02251_ _02252_ _02253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07592_ _02933_ _03012_ _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09400_ _03740_ ci_neuron.input_memory\[1\]\[4\] _00768_ _01874_ _04622_ _04623_
+ _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06543_ _02094_ _02142_ _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09331_ _04566_ _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_48_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06474_ _02117_ _00230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09262_ _04166_ _04138_ _04127_ _04536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05425_ ci_neuron.uut_simple_neuron.x2\[15\] _01096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08213_ ci_neuron.uut_simple_neuron.x0\[5\] _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09193_ _03967_ _04496_ _04497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05356_ _01027_ _01028_ _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08144_ _03680_ _03681_ _03683_ _03684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_114_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05287_ _00864_ _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08075_ _03606_ _03615_ _03626_ _03627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_31_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07026_ _02128_ _02603_ _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__04860__I _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09529__A2 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08977_ _04336_ _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07960__A1 _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07928_ _03504_ _00135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07859_ ci_neuron.uut_simple_neuron.titan_id_2\[6\] ci_neuron.uut_simple_neuron.titan_id_5\[6\]
+ _03447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_78_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09529_ _04724_ _04740_ _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08512__I0 _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09465__A1 ci_neuron.output_memory\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10235_ _00131_ net211 ci_neuron.uut_simple_neuron.titan_id_6\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10166_ _00092_ net210 ci_neuron.uut_simple_neuron.titan_id_2\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10097_ _00163_ net265 ci_neuron.uut_simple_neuron.titan_id_4\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_128_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04945__I _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06190_ _01820_ _01840_ _01841_ _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_79_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05210_ _00886_ _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05141_ _00743_ _00798_ _00820_ _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_4_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05072_ _00755_ _00160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09926__CLK net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08900_ _04293_ _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09880_ _00040_ net25 ci_neuron.value_i\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08831_ _04122_ ci_neuron.uut_simple_neuron.x2\[31\] _04210_ _04253_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07942__A1 _03512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05974_ _01601_ _01632_ _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08762_ _03955_ _04209_ _04213_ _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07713_ ci_neuron.uut_simple_neuron.titan_id_4\[12\] ci_neuron.uut_simple_neuron.titan_id_3\[12\]
+ _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08498__A2 _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08693_ internal_ih.spi_tx_byte_o\[3\] _04137_ _04157_ _04155_ _04158_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_04925_ _00639_ _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07644_ _03263_ _03266_ _03268_ _03269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08528__S _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04856_ _00597_ _00602_ _00606_ internal_ih.byte7\[0\] _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_0_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07575_ _02081_ _02480_ _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06526_ _02125_ _02128_ _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09314_ _04046_ ci_neuron.input_memory\[1\]\[16\] _04567_ _04569_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06457_ _01880_ _01963_ _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09245_ _04526_ _00469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05408_ _01038_ _01062_ _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06388_ _02030_ _02016_ _02032_ _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09176_ _04484_ _00442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05339_ _00812_ _00847_ _00867_ _01011_ _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_08127_ _03670_ _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08058_ _03611_ _03612_ _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07009_ _02519_ _02518_ _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_112_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10020_ ci_neuron.input_memory\[1\]\[20\] net109 ci_neuron.uut_simple_neuron.titan_id_1\[22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05475__A2 _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__04986__A1 internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10218_ _00115_ net241 ci_neuron.uut_simple_neuron.titan_id_5\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10149_ _00214_ net247 ci_neuron.uut_simple_neuron.titan_id_3\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09516__I2 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05690_ _01353_ _01354_ _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_89_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08575__C _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07360_ _02986_ _02987_ _02910_ _02978_ _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_45_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06311_ _01957_ _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07291_ _02897_ _02908_ _02919_ _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_115_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09030_ _04377_ _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06242_ _01825_ _01852_ _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_60_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06173_ _01825_ _01822_ _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05124_ _00786_ _00802_ _00803_ _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_13_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06966__A2 _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05055_ _00739_ _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09932_ _00447_ net170 ci_neuron.uut_simple_neuron.x0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08168__A1 _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09863_ _00442_ net69 ci_neuron.output_memory\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08814_ _04085_ _01433_ _04239_ _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_5_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09794_ _00373_ net53 internal_ih.byte5\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08745_ internal_ih.received_byte_count\[4\] _04199_ internal_ih.received_byte_count\[5\]
+ _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05957_ _01614_ _01615_ _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05888_ _01548_ _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08676_ internal_ih.spi_tx_byte_o\[0\] _04137_ _04142_ _04143_ _04144_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_04908_ _00642_ _00023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07627_ _03157_ _03193_ _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04839_ _00583_ internal_ih.received_byte_count\[2\] _00585_ _00590_ _00591_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07558_ _03182_ _03183_ _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06509_ _02130_ _02151_ _02152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07489_ _03109_ _03115_ _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_91_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07896__I _03478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08643__A2 _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09228_ _04059_ _03841_ _04514_ _04517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_121_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09159_ ci_neuron.uut_simple_neuron.titan_id_6\[23\] _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08520__I _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10003_ ci_neuron.input_memory\[1\]\[3\] net201 ci_neuron.uut_simple_neuron.titan_id_1\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_125_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05393__A1 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06645__A1 _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09673__D _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09526__I _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06860_ _02494_ _02495_ _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_87_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05811_ _01472_ _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_2_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06791_ _01983_ _02009_ _02428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05742_ _01405_ _00213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08530_ _04000_ _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_05673_ _01103_ _01332_ _01337_ _01338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08461_ _03735_ _03958_ _03959_ _03960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07412_ _02998_ _03039_ _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08392_ _03897_ _00187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07343_ _02962_ _02971_ _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07274_ _01920_ _02903_ _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06225_ _01872_ _01874_ _01875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_73_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09013_ _04357_ _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06156_ _01615_ _01766_ _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06087_ _01741_ _01742_ _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05107_ _00773_ _00757_ _00768_ _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09915_ _00011_ net16 ci_neuron.address_i\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05038_ _00722_ _00723_ _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09846_ _00425_ net208 ci_neuron.output_memory\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08561__A1 _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06989_ ci_neuron.uut_simple_neuron.x3\[21\] _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05375__A1 _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09777_ _00356_ net64 internal_ih.byte3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08728_ _04178_ net31 _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_107_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08659_ spi_interface_cvonk.state\[2\] spi_interface_cvonk.state\[1\] _04127_ _04128_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_37_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09655__I1 ci_neuron.output_memory\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06010_ _01667_ _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07043__A1 _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07961_ _03532_ _00141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06912_ _02500_ _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09700_ spi_interface_cvonk.SS_r\[1\] net121 spi_interface_cvonk.SS_r\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07892_ _03475_ _00128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06843_ _02477_ _02478_ _02479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09631_ _04813_ _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06774_ _02411_ _02356_ _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09562_ _03904_ ci_neuron.input_memory\[1\]\[28\] _01792_ _03230_ _04760_ _04761_
+ _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA_fanout52_I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08513_ _04004_ _00259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05725_ _01218_ _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05109__A1 _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09343__I0 _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07649__A3 _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09493_ _04697_ _04707_ _04709_ _04710_ _00533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05656_ _00888_ _01174_ _01320_ _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08444_ _03942_ _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05587_ _01212_ _01253_ _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08375_ _03881_ _03882_ _03883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07326_ _02332_ _02882_ _02955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09646__I1 ci_neuron.output_memory\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07257_ _01908_ _02828_ _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07188_ _02282_ _02818_ _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06208_ ci_neuron.uut_simple_neuron.x3\[3\] ci_neuron.uut_simple_neuron.x3\[4\] _01859_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_60_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06139_ _01792_ _01793_ _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05694__I _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05596__A1 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09829_ _00408_ net126 internal_ih.spi_tx_byte_o\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09334__I0 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout60 net61 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout71 net72 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09637__I1 ci_neuron.output_memory\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout82 net83 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout93 net94 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08773__A1 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09951__D _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09325__I0 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06490_ _02131_ _02132_ _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05510_ _00858_ _01178_ _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_75_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05441_ _01108_ _01111_ _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09628__I1 ci_neuron.output_memory\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08160_ _03692_ _03695_ _03696_ _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07111_ _02724_ _02742_ _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_82_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05372_ _01042_ _01019_ _01043_ _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08091_ _03639_ _03640_ _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07042_ _02672_ _02673_ _02674_ _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05814__A2 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07016__A1 _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08764__A1 _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08993_ internal_ih.current_instruction\[4\] _04340_ _04346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07944_ ci_neuron.uut_simple_neuron.titan_id_2\[20\] ci_neuron.uut_simple_neuron.titan_id_5\[20\]
+ _03518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07875_ _03453_ _03459_ _03460_ _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06826_ _02462_ _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09614_ _04803_ _00561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09316__I0 _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04858__I _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06757_ _02135_ _02394_ _02395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09545_ _04743_ _04751_ _04753_ _04754_ _00541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06688_ _02282_ _02326_ _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_104_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05708_ _01191_ _01335_ _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09476_ _04673_ _04690_ _04694_ _04695_ _00531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_109_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05639_ _01240_ _01278_ _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05502__A1 _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08427_ _03925_ _03926_ _03927_ _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_108_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08358_ _03862_ _03864_ _03867_ _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_19_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07309_ ci_neuron.uut_simple_neuron.x3\[25\] _02937_ _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08289_ _03807_ _00174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10251_ _00148_ net51 ci_neuron.uut_simple_neuron.titan_id_6\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10182_ _00080_ net99 ci_neuron.uut_simple_neuron.titan_id_2\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout250 net251 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout261 net263 net261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout283 net284 net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout272 net284 net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05990_ _01449_ _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09681__D _00268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04941_ internal_ih.byte6\[6\] _00658_ _00659_ internal_ih.byte2\[6\] _00662_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07660_ ci_neuron.uut_simple_neuron.titan_id_4\[3\] ci_neuron.uut_simple_neuron.titan_id_3\[3\]
+ _03282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_04872_ _00618_ _00029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07591_ _03148_ _03149_ _03212_ _03216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06611_ _02167_ _02207_ _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05732__A1 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06542_ _02045_ _02145_ _02183_ _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_75_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09330_ _04577_ _00503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09261_ _04534_ _04184_ _04124_ _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09474__A2 _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06473_ _02070_ _02116_ _02117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08212_ _03739_ _03740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05424_ _00860_ _01090_ _01094_ _01095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_7_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09192_ _04487_ _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05355_ _00993_ _00994_ _01026_ _01028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08143_ ci_neuron.uut_simple_neuron.titan_id_1\[23\] ci_neuron.uut_simple_neuron.titan_id_0\[23\]
+ _03683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_15_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08074_ _03614_ _03617_ _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08985__A1 _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07025_ _02606_ _02632_ _02657_ _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05286_ _00935_ _00946_ _00947_ _00949_ _00959_ _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09444__I _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08976_ internal_ih.byte7\[5\] internal_ih.byte6\[5\] _04332_ _04336_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07927_ _03502_ _03503_ _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07858_ _03442_ _03445_ _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07789_ _03389_ _00112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06809_ _02383_ _02445_ _02446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_97_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09528_ _03864_ ci_neuron.input_memory\[1\]\[23\] _01433_ _02928_ _04738_ _04739_
+ _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_39_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08512__I1 _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07476__A1 _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09459_ _04673_ _04676_ _04679_ _04681_ _00528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_93_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07139__I _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10234_ _00130_ net211 ci_neuron.uut_simple_neuron.titan_id_6\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10165_ _00091_ net209 ci_neuron.uut_simple_neuron.titan_id_2\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10096_ _00162_ net276 ci_neuron.uut_simple_neuron.titan_id_4\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_128_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09456__A2 _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05140_ _00735_ _00813_ _00816_ _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_52_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05071_ _00752_ _00754_ _00755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08830_ _04252_ _00328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05973_ _01604_ _01631_ _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08761_ _00745_ _04211_ _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07712_ _03322_ _03324_ _03325_ _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_79_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08692_ _04141_ _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04924_ _00651_ _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07643_ _03176_ _03179_ _03267_ _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04855_ _00605_ _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05705__B2 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07574_ _03198_ _03199_ _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08608__I _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09313_ _04568_ _00495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09447__A2 _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06525_ _02073_ _02159_ _02158_ _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__07458__A1 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06456_ _01876_ _02100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09244_ _04094_ _03893_ _04525_ _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05407_ _00959_ _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_60_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09175_ ci_neuron.uut_simple_neuron.titan_id_6\[31\] _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06387_ _02013_ _02031_ _02012_ _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08126_ _03668_ _03669_ _03670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05338_ _00983_ _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07630__A1 _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05269_ _00941_ _00943_ _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08057_ ci_neuron.uut_simple_neuron.titan_id_1\[9\] ci_neuron.uut_simple_neuron.titan_id_0\[9\]
+ _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07008_ _02576_ _02588_ _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_112_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07933__A2 ci_neuron.uut_simple_neuron.titan_id_5\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09174__I _04483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05944__A1 _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08959_ _04326_ _00383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09438__A2 _04662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10217_ _00114_ net237 ci_neuron.uut_simple_neuron.titan_id_5\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10148_ _00213_ net247 ci_neuron.uut_simple_neuron.titan_id_3\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10079_ _00176_ net113 ci_neuron.uut_simple_neuron.titan_id_0\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09516__I3 _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07290_ _02852_ _02896_ _02919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06310_ _01868_ _01934_ _01956_ _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06241_ _01889_ _01863_ _01885_ _01890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_127_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05787__I _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06172_ ci_neuron.uut_simple_neuron.x3\[0\] _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05123_ _00789_ _00799_ _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_123_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05054_ _00738_ _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09931_ _00446_ net170 ci_neuron.uut_simple_neuron.x0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09862_ _00441_ net69 ci_neuron.output_memory\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08813_ _04079_ _04211_ _04243_ _00320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09793_ _00372_ net55 internal_ih.byte5\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05956_ _01327_ _01478_ _01524_ _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_08744_ _04194_ _04200_ _00294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08539__S _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04907_ internal_ih.byte5\[0\] _00640_ _00641_ internal_ih.byte1\[0\] _00642_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05887_ _01511_ _01512_ _01546_ _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08675_ internal_ih.spi_rx_byte_i\[0\] _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07626_ _03249_ _03250_ _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04838_ _00586_ _00588_ _00589_ _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07557_ _02082_ _03113_ _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06508_ _02134_ _02150_ _02151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_75_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07488_ _03112_ _03114_ _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06439_ _02081_ _02082_ _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09227_ _04516_ _00461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09158_ _04475_ _00433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08109_ _03655_ _00072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08651__I0 ci_neuron.uut_simple_neuron.x0\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09089_ ci_neuron.output_val_internal\[29\] ci_neuron.output_val_internal\[21\] ci_neuron.output_val_internal\[13\]
+ ci_neuron.output_val_internal\[5\] _04366_ _04367_ _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_101_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08801__I _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10002_ ci_neuron.input_memory\[1\]\[2\] net200 ci_neuron.uut_simple_neuron.titan_id_1\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_125_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_26_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08945__I1 internal_ih.byte4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05810_ ci_neuron.uut_simple_neuron.x2\[24\] _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06790_ _02425_ _02426_ _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05741_ _01400_ _01404_ _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05672_ _01336_ _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08460_ _03942_ _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07411_ _03028_ _03038_ _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_35_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08391_ _03890_ _03892_ _03896_ _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07342_ _02963_ _02970_ _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07273_ _01895_ _01899_ _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_98_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06224_ _01873_ _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09012_ internal_ih.data_pointer\[0\] _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06155_ _01613_ _01765_ _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05106_ _00781_ _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_44_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06086_ _01412_ _01697_ _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09914_ _00010_ net13 ci_neuron.address_i\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05037_ ci_neuron.address_i\[1\] ci_neuron.address_i\[0\] ci_neuron.address_i\[2\]
+ _00723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09845_ _00424_ net208 ci_neuron.output_memory\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06988_ _02616_ _02556_ _02621_ _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09776_ _00355_ net50 internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05939_ _01597_ _01598_ _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_68_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08727_ _04177_ _04186_ _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_107_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08313__A2 _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_53_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08658_ spi_interface_cvonk.state\[0\] _04127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_37_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ _03168_ _03169_ _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_120_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08589_ _04011_ _04069_ _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__04886__A1 internal_ih.byte4\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04886__B2 internal_ih.byte0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_62_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09362__I _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06315__A1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__04877__B2 _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07960_ _03530_ _03531_ _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06911_ _02505_ _02508_ _02545_ _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07891_ _03473_ _03474_ _03475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06842_ _02040_ _02437_ _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09272__I _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09630_ ci_neuron.stream_o\[17\] ci_neuron.output_memory\[17\] _04811_ _04813_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06773_ _02355_ _02411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09561_ _04700_ _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05724_ _01369_ _01387_ _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08512_ _04003_ _02089_ _03969_ _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09343__I1 ci_neuron.input_memory\[1\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06306__A1 _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09492_ ci_neuron.output_val_internal\[17\] _04705_ _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05655_ _01083_ _01210_ _01176_ _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_34_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08443_ _03943_ _03944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_05586_ _00860_ _01207_ _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08374_ _03869_ _03872_ _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07325_ _02341_ _02881_ _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08854__I0 internal_ih.byte1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07256_ _02273_ _02291_ _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06207_ _01821_ _01843_ _01839_ _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_5_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07187_ _02288_ _02817_ _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06580__B _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07034__A2 _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06138_ ci_neuron.uut_simple_neuron.x2\[30\] _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06069_ _01594_ _01725_ _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05596__A2 _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09761__CLK net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09828_ _00407_ net139 internal_ih.spi_tx_byte_o\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09759_ _00338_ net67 internal_ih.byte1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_68_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08845__I0 internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout61 net62 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout50 net51 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout72 net73 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout83 net84 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_70_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xfanout94 net96 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05339__A2 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07605__I ci_neuron.uut_simple_neuron.x3\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05440_ _01109_ _01110_ _01061_ _01059_ _01008_ _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_129_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05371_ _01002_ _01011_ _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07110_ _02739_ _02741_ _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05275__A1 _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08090_ ci_neuron.uut_simple_neuron.titan_id_1\[14\] ci_neuron.uut_simple_neuron.titan_id_0\[14\]
+ _03640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07041_ _02619_ _02627_ _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__04873__I1 internal_ih.byte3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08992_ _04345_ _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07943_ _03515_ _03516_ _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06527__A1 _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07874_ ci_neuron.uut_simple_neuron.titan_id_2\[7\] ci_neuron.uut_simple_neuron.titan_id_5\[7\]
+ ci_neuron.uut_simple_neuron.titan_id_2\[6\] ci_neuron.uut_simple_neuron.titan_id_5\[6\]
+ _03460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_06825_ _02418_ _02461_ _02462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09613_ ci_neuron.stream_o\[10\] ci_neuron.output_memory\[10\] _04800_ _04803_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06756_ _02096_ _02230_ _02394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_09544_ ci_neuron.output_val_internal\[25\] _04749_ _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06687_ _02182_ _02287_ _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05707_ _01188_ _01370_ _01104_ _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_66_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09475_ ci_neuron.output_val_internal\[15\] _04680_ _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05638_ _01300_ _01303_ _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_65_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08426_ _00709_ _03923_ _00728_ _00714_ _03927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_05569_ _01169_ _01197_ _01237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08827__I0 _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08357_ _03865_ _03866_ _03867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07308_ ci_neuron.uut_simple_neuron.x3\[26\] _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08288_ _03803_ _03806_ _03807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07239_ ci_neuron.uut_simple_neuron.x3\[24\] _02868_ _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10250_ _00147_ net80 ci_neuron.uut_simple_neuron.titan_id_6\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09252__I0 _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10181_ _00079_ net99 ci_neuron.uut_simple_neuron.titan_id_2\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout240 net241 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout251 net252 net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout262 net263 net262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout273 net275 net273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout284 net285 net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07191__A1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04940_ _00661_ _00014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_04871_ internal_ih.byte7\[4\] _00616_ _00617_ _00610_ _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07590_ _03215_ _00248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06610_ _02167_ _02207_ _02251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06541_ _02181_ _02182_ _02183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_9_Left_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06472_ _02072_ _02115_ _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_62_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09260_ spi_interface_cvonk.SS_r\[2\] _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_117_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05423_ _01018_ _01093_ _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08211_ ci_neuron.uut_simple_neuron.x0\[4\] _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08682__A1 _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09191_ _03961_ _04494_ _04495_ _00446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05354_ _00993_ _00994_ _01026_ _01027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_16_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08142_ _03682_ _00079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05285_ _00879_ _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08073_ _03625_ _00095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07024_ _02608_ _02631_ _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06748__A1 _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08975_ _04335_ _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07926_ ci_neuron.uut_simple_neuron.titan_id_2\[17\] ci_neuron.uut_simple_neuron.titan_id_5\[17\]
+ _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07857_ _03443_ _03444_ _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07788_ _03387_ _03388_ _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06808_ _02388_ _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_97_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06739_ _02332_ _02341_ _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09527_ _04668_ _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_42_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09458_ ci_neuron.output_val_internal\[12\] _04680_ _04681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09389_ ci_neuron.output_memory\[3\] _04600_ _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08409_ ci_neuron.uut_simple_neuron.x0\[28\] ci_neuron.uut_simple_neuron.x0\[29\]
+ _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_22_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06739__A1 _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08728__A2 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10233_ _00129_ net193 ci_neuron.uut_simple_neuron.titan_id_6\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10164_ _00090_ net209 ci_neuron.uut_simple_neuron.titan_id_2\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10095_ ci_neuron.uut_simple_neuron.x3\[0\] net264 ci_neuron.uut_simple_neuron.titan_id_4\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_128_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09370__I _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06978__A1 _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05070_ _00733_ _00753_ _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05972_ _01607_ _01630_ _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08760_ _03947_ _04209_ _04212_ _00298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07155__A1 _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07711_ ci_neuron.uut_simple_neuron.titan_id_4\[11\] ci_neuron.uut_simple_neuron.titan_id_3\[11\]
+ _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08691_ _04134_ _04154_ _04156_ _00285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04923_ internal_ih.byte5\[7\] _00646_ _00647_ internal_ih.byte1\[7\] _00651_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07642_ _03162_ _03174_ _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04854_ _00604_ _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07573_ _03109_ _03115_ _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09312_ _04040_ ci_neuron.input_memory\[1\]\[15\] _04567_ _04568_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06524_ _02119_ _02163_ _02165_ _02166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07458__A2 _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05469__A1 _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06455_ _02088_ _02098_ _02099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_75_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09243_ _04487_ _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06386_ _01947_ _01971_ _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05406_ _01076_ _01064_ _01077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09174_ _04483_ _00441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05337_ _01006_ _01008_ _01009_ _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08125_ ci_neuron.uut_simple_neuron.titan_id_1\[20\] ci_neuron.uut_simple_neuron.titan_id_0\[20\]
+ _03669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_16_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05268_ _00909_ _00942_ _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08056_ _03609_ _03610_ _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07007_ _02637_ _02640_ _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_113_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05199_ _00876_ _00226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_112_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08430__I1 _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08958_ internal_ih.byte6\[5\] internal_ih.byte5\[5\] _04322_ _04326_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07909_ _03485_ _03487_ _03488_ _03489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08889_ internal_ih.byte2\[7\] internal_ih.byte1\[7\] _04285_ _04287_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09446__I0 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09461__I3 _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06989__I ci_neuron.uut_simple_neuron.x3\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10216_ _00113_ net236 ci_neuron.uut_simple_neuron.titan_id_5\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09365__I _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10147_ _00212_ net245 ci_neuron.uut_simple_neuron.titan_id_3\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_7_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10078_ _00175_ net173 ci_neuron.uut_simple_neuron.titan_id_0\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06360__A2 _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_99_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06240_ _01857_ _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_73_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06171_ _01824_ _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07612__A2 _03233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05122_ _00789_ _00799_ _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05053_ ci_neuron.uut_simple_neuron.x2\[1\] _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05623__A1 _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09930_ _00445_ net189 ci_neuron.uut_simple_neuron.x0\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09861_ _00440_ net80 ci_neuron.output_memory\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08812_ _01381_ _04221_ _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09792_ _00371_ net41 internal_ih.byte5\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05955_ _01580_ _01613_ _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08743_ internal_ih.received_byte_count\[4\] _04199_ _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_04906_ _00627_ _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05886_ _01511_ _01512_ _01546_ _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08674_ _04141_ _04142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07625_ _02121_ _03204_ _03250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04837_ internal_ih.expected_byte_count\[3\] _00584_ internal_ih.received_byte_count\[5\]
+ internal_ih.received_byte_count\[1\] _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07556_ _02489_ _02507_ _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06507_ _02147_ _02149_ _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07487_ _02082_ _03113_ _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07300__A1 _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09226_ _04052_ _03840_ _04514_ _04516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06438_ _02053_ _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07851__A2 ci_neuron.uut_simple_neuron.titan_id_5\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06369_ _02012_ _02014_ _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09157_ ci_neuron.uut_simple_neuron.titan_id_6\[22\] _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08108_ _03652_ _03654_ _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09088_ _04417_ ci_neuron.stream_o\[5\] ci_neuron.stream_o\[21\] _04418_ _04430_
+ _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_32_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08039_ ci_neuron.uut_simple_neuron.titan_id_1\[6\] ci_neuron.uut_simple_neuron.titan_id_0\[6\]
+ _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10001_ ci_neuron.input_memory\[1\]\[1\] net200 ci_neuron.uut_simple_neuron.titan_id_1\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_125_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05740_ _01313_ _01401_ _01403_ _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08439__I _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05671_ _01333_ _01335_ _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07410_ _03031_ _03037_ _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08390_ _03894_ _03895_ _03896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07341_ _02966_ _02969_ _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_73_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07272_ _02900_ _02901_ _02902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06223_ ci_neuron.uut_simple_neuron.x3\[4\] _01873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09011_ internal_ih.data_pointer\[1\] internal_ih.data_pointer\[0\] _04359_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06154_ _01756_ _01759_ _01808_ _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05105_ _00779_ _00785_ _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06085_ _01557_ _01696_ _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09913_ _00009_ net6 ci_neuron.address_i\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05036_ ci_neuron.address_i\[22\] ci_neuron.address_i\[23\] _00716_ _00721_ _00722_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09844_ _00423_ net195 ci_neuron.output_memory\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06987_ _02551_ _02620_ _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09775_ _00354_ net50 internal_ih.byte3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05938_ _01547_ _01552_ _01548_ _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08726_ _04178_ _04183_ _04185_ _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_107_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05869_ _01529_ _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08657_ spi_interface_cvonk.SCLK_r\[2\] _04125_ _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07608_ _03231_ _03232_ _03233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08588_ _03996_ _04067_ _04068_ _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_48_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07539_ _03163_ _03164_ _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09209_ _04506_ _00453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_106_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07856__C ci_neuron.uut_simple_neuron.titan_id_5\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06315__A2 _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06910_ _02497_ _02504_ _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07890_ ci_neuron.uut_simple_neuron.titan_id_2\[10\] ci_neuron.uut_simple_neuron.titan_id_5\[10\]
+ _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09553__I _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06841_ _02041_ _02436_ _02477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06772_ _02406_ _02409_ _02410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09560_ ci_neuron.output_memory\[28\] _04766_ _04767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05723_ _01374_ _01378_ _01386_ _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09491_ _04701_ _04708_ _04709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08511_ _03996_ _03998_ _03999_ _04002_ _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XANTENNA__07503__A1 _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08442_ _03942_ _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05654_ _01318_ _01296_ _01297_ _01284_ _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA_fanout38_I ci_neuron.uut_simple_neuron.x2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05585_ _01179_ _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08373_ _03863_ _03874_ _03881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07324_ _02951_ _02952_ _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07255_ _02855_ _02884_ _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_61_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08854__I1 internal_ih.byte0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06206_ _01856_ _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07186_ _02441_ _02740_ _02816_ _02817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_42_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06137_ _01668_ _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_57_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06068_ _01691_ _01724_ _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05019_ ci_neuron.uut_simple_neuron.x0\[1\] _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09827_ _00406_ net125 internal_ih.spi_tx_byte_o\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08790__I0 _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09758_ _00337_ net123 internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08709_ _04167_ _04169_ _04130_ _00290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09689_ _00276_ net221 ci_neuron.uut_simple_neuron.x3\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_68_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout40 net42 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout62 net72 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout51 net52 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout73 net119 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout95 net96 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout84 net97 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout242_I net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09238__A1 _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05370_ _01039_ _01040_ _01041_ _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_16_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07040_ _02629_ _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09410__A1 ci_neuron.output_memory\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08991_ _04155_ internal_ih.current_instruction\[3\] _04339_ _04345_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07942_ _03512_ _03513_ _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07873_ _03457_ _03458_ _03459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06824_ _02422_ _02460_ _02461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09612_ _04802_ _00560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09543_ _04746_ _04752_ _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06755_ _02382_ _02392_ _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_92_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06686_ _01928_ _02324_ _02325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_104_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05706_ _01191_ _01335_ _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_09474_ _04677_ _04693_ _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_47_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05637_ _01078_ _01301_ _01302_ _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08425_ _00708_ _00709_ ci_neuron.stream_enabled _03923_ _03926_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_108_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08356_ _03856_ _03859_ _03866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07307_ _02928_ _02869_ _02935_ _02936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05568_ _00959_ _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08827__I1 _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05499_ _01134_ _01155_ _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08287_ _03804_ _03805_ _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_6_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07238_ ci_neuron.uut_simple_neuron.x3\[25\] _02868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07169_ ci_neuron.uut_simple_neuron.x3\[23\] ci_neuron.uut_simple_neuron.x3\[24\]
+ _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_61_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09252__I1 _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07963__A1 _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10180_ _00078_ net99 ci_neuron.uut_simple_neuron.titan_id_2\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout241 net242 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout230 net231 net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout252 net290 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout263 net285 net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout274 net275 net274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout285 net289 net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_57_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09368__I _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04870_ internal_ih.byte4\[4\] internal_ih.byte3\[4\] _00608_ _00617_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08648__S _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06540_ _02144_ _02182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06471_ _02112_ _02114_ _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05422_ _00982_ _01092_ _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08210_ _03738_ _00194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09190_ _03724_ _04491_ _04495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05353_ _00996_ _01025_ _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08141_ _03680_ _03681_ _03682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_125_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05284_ _00953_ _00956_ _00951_ _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08072_ _03623_ _03624_ _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07023_ _01857_ _02655_ _02656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08974_ internal_ih.byte7\[4\] internal_ih.byte6\[4\] _04332_ _04335_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06430__I _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07925_ _03500_ _03501_ _03502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07856_ ci_neuron.uut_simple_neuron.titan_id_2\[5\] ci_neuron.uut_simple_neuron.titan_id_5\[5\]
+ ci_neuron.uut_simple_neuron.titan_id_2\[4\] ci_neuron.uut_simple_neuron.titan_id_5\[4\]
+ _03444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07787_ ci_neuron.uut_simple_neuron.titan_id_4\[25\] ci_neuron.uut_simple_neuron.titan_id_3\[25\]
+ _03388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_06807_ _02280_ _02391_ _02443_ _02444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_97_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04999_ internal_ih.byte2\[7\] _00691_ _00695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06738_ _01958_ _02375_ _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_119_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09526_ _04666_ _04738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09457_ _04610_ _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_42_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06669_ _02301_ _02307_ _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_109_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08408_ _03903_ _03905_ _03911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09388_ _04598_ _04617_ _04619_ _04620_ _00518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_117_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08339_ _03850_ _03851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_22_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08092__I _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_128_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06987__A2 _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06739__A2 _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10232_ _00128_ net208 ci_neuron.uut_simple_neuron.titan_id_6\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10163_ _00089_ net209 ci_neuron.uut_simple_neuron.titan_id_2\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10094_ _00192_ net74 ci_neuron.uut_simple_neuron.titan_id_0\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_128_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06978__A2 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05971_ _01567_ _01629_ _01630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07710_ ci_neuron.uut_simple_neuron.titan_id_4\[11\] ci_neuron.uut_simple_neuron.titan_id_3\[11\]
+ _03324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10131__CLK net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08690_ _04155_ _04149_ _04156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04922_ _00650_ _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07641_ _03264_ _03189_ _03265_ _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04853_ _00594_ _00603_ _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07572_ _03112_ _03114_ _03198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06523_ _02120_ _02162_ _02165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09311_ _04566_ _04567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__04913__B2 internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06454_ _01966_ _02097_ _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09242_ _04524_ _00468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08905__I _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06385_ _02018_ _02019_ _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05405_ _01075_ _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09173_ ci_neuron.uut_simple_neuron.titan_id_6\[30\] _04483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05336_ _00852_ _00972_ _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08124_ ci_neuron.uut_simple_neuron.titan_id_1\[19\] ci_neuron.uut_simple_neuron.titan_id_0\[19\]
+ _03657_ _03665_ _03667_ _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_43_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05267_ _00914_ _00942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08055_ _03606_ _03607_ _03610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07006_ _02638_ _02573_ _02639_ _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05198_ _00851_ _00875_ _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_112_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08957_ _04325_ _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07908_ ci_neuron.uut_simple_neuron.titan_id_2\[13\] ci_neuron.uut_simple_neuron.titan_id_5\[13\]
+ _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09471__I _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08888_ _04286_ _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07146__A2 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07839_ ci_neuron.uut_simple_neuron.titan_id_2\[3\] ci_neuron.uut_simple_neuron.titan_id_5\[3\]
+ _03429_ _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_98_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08087__I _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09509_ _04700_ _04724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10215_ _00112_ net240 ci_neuron.uut_simple_neuron.titan_id_5\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07166__I ci_neuron.uut_simple_neuron.x3\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10146_ _00211_ net244 ci_neuron.uut_simple_neuron.titan_id_3\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05396__A1 _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10077_ _00174_ net173 ci_neuron.uut_simple_neuron.titan_id_0\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout155_I net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06170_ _01823_ _01824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_108_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05121_ _00801_ _00223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05052_ _00736_ _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09860_ _00439_ net81 ci_neuron.output_memory\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05387__A1 _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08811_ _04242_ _00319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09791_ _00370_ net43 internal_ih.byte5\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05954_ _01326_ _01612_ _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08742_ _04193_ _04198_ _04199_ _00293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08673_ _04138_ _04140_ _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_04905_ _00639_ _00640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout68_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07624_ _02131_ _02103_ _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05885_ _01076_ _01545_ _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_95_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04836_ internal_ih.expected_byte_count\[0\] _00587_ _00588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07555_ _03159_ _03180_ _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07486_ _02489_ _02507_ _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06506_ _01925_ _02148_ _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06437_ _02047_ _02081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07300__A2 _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09225_ _04515_ _00460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06368_ _01947_ _01971_ _02013_ _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09156_ _04474_ _00432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06299_ _01867_ _01936_ _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05319_ _00992_ _00203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08107_ _03653_ _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09087_ _04405_ _04429_ _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08038_ _03595_ _00090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_73_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09600__I1 ci_neuron.output_memory\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10000_ ci_neuron.input_memory\[1\]\[0\] net188 ci_neuron.uut_simple_neuron.titan_id_1\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09989_ _00504_ net91 ci_neuron.input_memory\[1\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06802__A1 _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10129_ _00161_ net265 ci_neuron.uut_simple_neuron.titan_id_3\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout272_I net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06869__A1 _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05670_ _01226_ _01290_ _01334_ _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07340_ _02967_ _02968_ _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07271_ _02824_ _02830_ _02901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09010_ _04357_ _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06222_ _01838_ _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06153_ _01714_ _01760_ _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05104_ _00780_ _00754_ _00782_ _00784_ _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_123_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06084_ _01738_ _01739_ _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05319__I _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09912_ _00008_ net6 ci_neuron.address_i\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05035_ _00717_ _00718_ _00719_ _00720_ _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_09843_ _00422_ net161 ci_neuron.output_memory\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06986_ _02555_ _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09774_ _00353_ net49 internal_ih.byte2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05937_ _01593_ _01596_ _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_69_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08725_ _04184_ _04140_ _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05868_ _01479_ _01525_ _01529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08656_ spi_interface_cvonk.SCLK_r\[1\] _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_107_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07607_ _03229_ _03230_ ci_neuron.uut_simple_neuron.x3\[29\] _03232_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08587_ ci_neuron.value_i\[20\] _04055_ _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_120_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07538_ _02870_ _03091_ _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05799_ _01377_ _01371_ _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07469_ _03094_ _03095_ _03096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09208_ _04003_ _03772_ _04488_ _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_121_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09139_ ci_neuron.uut_simple_neuron.titan_id_6\[13\] _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08785__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09585__I0 _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08776__A1 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout118_I net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10192__D _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07200__A1 _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06840_ _01847_ _02428_ _02475_ _02476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06771_ _02309_ _02407_ _02408_ _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05762__A1 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05722_ _01384_ _01385_ _01386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09490_ _03824_ ci_neuron.input_memory\[1\]\[17\] _01184_ _02445_ _04691_ _04692_
+ _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08510_ ci_neuron.value_i\[9\] _04001_ _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05653_ _01286_ _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08441_ _03925_ _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05584_ _01215_ _01249_ _01250_ _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_86_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08372_ _03876_ _03879_ _03880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07323_ _01948_ _02892_ _02952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07254_ _02879_ _02883_ _02884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_102_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06205_ _01852_ _01854_ _01855_ _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_60_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04876__I0 internal_ih.byte4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07185_ _02442_ _02615_ _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06136_ _01789_ _01767_ _01790_ _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_57_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06067_ _01650_ _01723_ _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05018_ _00705_ _00057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08519__A1 ci_neuron.value_i\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09826_ _00405_ net132 internal_ih.spi_tx_byte_o\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06969_ _02173_ _02148_ _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09757_ _00336_ net124 internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08708_ spi_interface_cvonk.buffer\[7\] _04168_ _04131_ _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09688_ _00275_ net221 ci_neuron.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05505__A1 _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08639_ _04110_ _03230_ _04111_ _04112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_81_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout30 net31 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout41 net42 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout63 net66 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout52 net73 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout74 net79 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout96 net97 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout85 net87 net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_92_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09573__I3 ci_neuron.uut_simple_neuron.x3\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05744__A1 _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05339__A4 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05027__A3 _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08990_ _04170_ _04340_ _04344_ _00396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07972__A2 ci_neuron.uut_simple_neuron.titan_id_5\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07941_ ci_neuron.uut_simple_neuron.titan_id_2\[19\] ci_neuron.uut_simple_neuron.titan_id_5\[19\]
+ _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07872_ _03447_ _03451_ _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06823_ _02424_ _02459_ _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09611_ ci_neuron.stream_o\[9\] ci_neuron.output_memory\[9\] _04800_ _04802_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06754_ _02280_ _02391_ _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09542_ _03893_ ci_neuron.input_memory\[1\]\[25\] _01573_ _02934_ _04738_ _04739_
+ _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_78_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05705_ _01341_ _01346_ _01367_ _01368_ _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_06685_ _01935_ _02323_ _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_104_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09473_ _03825_ ci_neuron.input_memory\[1\]\[15\] _01098_ _02387_ _04691_ _04692_
+ _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_59_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05636_ _01251_ _01275_ _01302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08424_ _00724_ _03924_ _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05567_ _01067_ _01234_ _01235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10097__D _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08355_ _03850_ ci_neuron.uut_simple_neuron.x0\[22\] _03865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07306_ _02863_ _02934_ _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_63_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05498_ _01134_ _01155_ _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08286_ _03783_ _03796_ _03794_ _03805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_116_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07237_ _02731_ _02864_ _02866_ _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07168_ _02734_ _02735_ _02798_ _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06119_ _01771_ _01774_ _01775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07099_ _02730_ _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout231 net233 net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout220 net225 net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout242 net251 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout253 net258 net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout264 net266 net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout286 net288 net286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout275 net276 net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09809_ _00388_ net54 internal_ih.byte7\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08818__I _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06390__A1 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06470_ _02113_ _02063_ _02114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_44_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05421_ _00964_ _01055_ _01091_ _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08140_ ci_neuron.uut_simple_neuron.titan_id_1\[23\] ci_neuron.uut_simple_neuron.titan_id_0\[23\]
+ _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05352_ _00905_ _01024_ _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05283_ _00957_ _00202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08071_ ci_neuron.uut_simple_neuron.titan_id_1\[11\] ci_neuron.uut_simple_neuron.titan_id_0\[11\]
+ _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07022_ _02653_ _02654_ _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08973_ _04334_ _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07924_ _03497_ _03498_ _03501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07855_ ci_neuron.uut_simple_neuron.titan_id_2\[5\] ci_neuron.uut_simple_neuron.titan_id_5\[5\]
+ _03443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07786_ ci_neuron.uut_simple_neuron.titan_id_4\[24\] ci_neuron.uut_simple_neuron.titan_id_3\[24\]
+ _03376_ _03384_ _03386_ _03387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_06806_ _02441_ _02442_ _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05184__A2 _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08638__I _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04998_ _00694_ _00047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06737_ _01968_ _02374_ _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_65_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09525_ ci_neuron.output_memory\[23\] _04722_ _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06668_ _02250_ _02253_ _02302_ _02304_ _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_66_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09456_ _04677_ _04678_ _04679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_109_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05619_ _01262_ _01271_ _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08407_ _03905_ ci_neuron.uut_simple_neuron.x0\[30\] _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06599_ _02219_ _02221_ _02239_ _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09387_ ci_neuron.output_val_internal\[2\] _04611_ _04620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08338_ ci_neuron.uut_simple_neuron.x0\[21\] _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_22_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07633__A1 _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08269_ _03782_ _03784_ _03778_ _03779_ _03777_ _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10231_ _00158_ net192 ci_neuron.uut_simple_neuron.titan_id_6\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07936__A2 ci_neuron.uut_simple_neuron.titan_id_5\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10162_ _00088_ net197 ci_neuron.uut_simple_neuron.titan_id_2\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10093_ _00191_ net74 ci_neuron.uut_simple_neuron.titan_id_0\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09528__I3 _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05970_ _01628_ _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04921_ internal_ih.byte5\[6\] _00646_ _00647_ internal_ih.byte1\[6\] _00650_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_49_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07640_ _03184_ _03191_ _03265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04852_ _00599_ _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07571_ _03195_ _03196_ _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06522_ _02164_ _00231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09310_ _04542_ _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06453_ _02093_ _02096_ _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09241_ _04089_ _03877_ _04519_ _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_113_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06384_ _01945_ _02021_ _02028_ _02015_ _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_91_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05404_ _01067_ _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09172_ _04482_ _00440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07615__A1 _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05335_ _00964_ _01007_ _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_60_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08123_ _03660_ _03666_ _03667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08054_ ci_neuron.uut_simple_neuron.titan_id_1\[8\] ci_neuron.uut_simple_neuron.titan_id_0\[8\]
+ _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07005_ _02569_ _02572_ _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05266_ _00938_ _00940_ _00941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05197_ _00854_ _00874_ _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_112_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08956_ internal_ih.byte6\[4\] internal_ih.byte5\[4\] _04322_ _04325_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07907_ ci_neuron.uut_simple_neuron.titan_id_2\[13\] ci_neuron.uut_simple_neuron.titan_id_5\[13\]
+ _03487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08887_ internal_ih.byte2\[6\] internal_ih.byte1\[6\] _04285_ _04286_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06354__A1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07838_ _03425_ _03427_ _03428_ _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_27_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07769_ ci_neuron.uut_simple_neuron.titan_id_4\[22\] ci_neuron.uut_simple_neuron.titan_id_3\[22\]
+ _03372_ _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_27_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09508_ ci_neuron.output_memory\[20\] _04722_ _04723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_123_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09439_ ci_neuron.output_val_internal\[10\] _04655_ _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10214_ _00111_ net247 ci_neuron.uut_simple_neuron.titan_id_5\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10145_ _00210_ net243 ci_neuron.uut_simple_neuron.titan_id_3\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10076_ _00173_ net176 ci_neuron.uut_simple_neuron.titan_id_0\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08893__I0 internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05120_ _00778_ _00800_ _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08645__I0 _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05051_ _00735_ _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07357__I _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08810_ _04074_ _01368_ _04239_ _04242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08573__A2 _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09790_ _00369_ net43 internal_ih.byte4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05953_ ci_neuron.uut_simple_neuron.x2\[23\] _01379_ _01524_ _01612_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08741_ internal_ih.received_byte_count\[3\] _04197_ _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05884_ _01515_ _01544_ _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_84_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04904_ _00604_ _00639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08672_ spi_interface_cvonk.state\[2\] _04139_ _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07623_ _03246_ _03247_ _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04835_ internal_ih.received_byte_count\[0\] _00587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07554_ _03176_ _03179_ _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04898__B2 internal_ih.byte0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07485_ _03110_ _03111_ _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06505_ _01905_ _02000_ _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_52_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06436_ _01833_ _02079_ _02080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_91_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09224_ _04046_ _03822_ _04514_ _04515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06367_ _01951_ _01970_ _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09155_ ci_neuron.uut_simple_neuron.titan_id_6\[21\] _04474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06298_ _01944_ _01940_ _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05318_ _00958_ _00991_ _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08106_ ci_neuron.uut_simple_neuron.titan_id_1\[17\] ci_neuron.uut_simple_neuron.titan_id_0\[17\]
+ _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09086_ _04419_ ci_neuron.stream_o\[13\] _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05249_ _00885_ _00923_ _00924_ _00901_ _00855_ _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_08037_ _03593_ _03594_ _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09988_ _00503_ net92 ci_neuron.input_memory\[1\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08939_ _04315_ _00374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08098__I _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08875__I0 internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10128_ _00160_ net265 ci_neuron.uut_simple_neuron.titan_id_3\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10059_ _00544_ net103 ci_neuron.output_val_internal\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06869__A2 _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout265_I net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05541__A2 _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08866__I0 internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07270_ _02827_ _02829_ _02900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06221_ _01870_ _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06152_ _01648_ _01806_ _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08471__I _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06083_ _01604_ _01723_ _01739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05103_ _00783_ _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09911_ _00007_ net7 ci_neuron.address_i\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05034_ ci_neuron.address_i\[9\] ci_neuron.address_i\[8\] ci_neuron.address_i\[7\]
+ ci_neuron.address_i\[6\] _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_41_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09842_ _00421_ net192 ci_neuron.output_memory\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_13_Left_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09773_ _00352_ net48 internal_ih.byte2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06985_ _02442_ _02558_ _02618_ _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08724_ spi_interface_cvonk.SCLK_r\[2\] _04125_ _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05936_ _01594_ _01545_ _01595_ _01596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05867_ _01477_ _01479_ _01480_ _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08655_ spi_interface_cvonk.SS_r\[1\] _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07606_ _03229_ _03230_ _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08586_ _03848_ _04066_ _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_37_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07537_ _03087_ _03089_ _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05798_ _01458_ _01459_ _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07468_ _02682_ _02930_ _03095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08482__A1 _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07399_ _03004_ _03021_ _03026_ _03027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06419_ _02029_ _02033_ _02063_ _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_91_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09207_ _03994_ _04503_ _04505_ _00452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09138_ _04465_ _00423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09477__I _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09069_ internal_ih.spi_tx_byte_o\[3\] _04379_ _04414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06260__A3 _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_31_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05220__A1 _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08556__I _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_40_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06770_ _02351_ _02353_ _02408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05721_ _00740_ _01343_ _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05652_ _01075_ _01299_ _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08440_ _03940_ _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_81_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05583_ _01217_ _01231_ _01250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08371_ _03878_ _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07322_ _02323_ _02344_ _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07253_ _02332_ _02882_ _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_121_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07184_ _02796_ _02811_ _02814_ _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_104_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06204_ _01825_ _01845_ _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_60_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06135_ _01753_ _01761_ _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_57_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06066_ _01694_ _01722_ _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05017_ internal_ih.byte3\[7\] _00701_ _00705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08519__A2 _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09825_ _00404_ net131 internal_ih.spi_tx_byte_o\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06968_ _02600_ _02601_ _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09756_ _00335_ net123 internal_ih.byte0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09687_ _00274_ net221 ci_neuron.uut_simple_neuron.x3\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05919_ ci_neuron.uut_simple_neuron.x2\[26\] _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08707_ _04166_ _04141_ _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06899_ _02532_ _02533_ _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ _03939_ _04111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_83_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08569_ _03968_ _04053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_65_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout31 net35 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout20 net22 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout53 net55 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout42 net43 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout64 net66 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout97 net118 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout86 net88 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout75 net79 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_122_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08446__A1 ci_neuron.value_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09246__I0 _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05680__A1 _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05432__A1 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07940_ _03514_ _00137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07871_ _03455_ _03456_ _03445_ _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06822_ _02431_ _02458_ _02459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09610_ _04801_ _00559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06753_ _02386_ _02390_ _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09541_ ci_neuron.output_memory\[25\] _04744_ _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05704_ _01344_ _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_104_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06684_ _02044_ _02290_ _02322_ _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_78_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09472_ _04668_ _04692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout43_I net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05635_ _01251_ _01275_ _01301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08423_ _00714_ _03923_ _00710_ _03924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05566_ _01206_ _01233_ _01234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08354_ _03863_ _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07305_ _02868_ _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_63_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05497_ _01164_ _01165_ _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08285_ _03794_ ci_neuron.uut_simple_neuron.x0\[13\] _03790_ _03791_ _03789_ _03804_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_46_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07236_ _02797_ _02865_ _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_61_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07167_ _02730_ _02797_ _02798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_42_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06118_ _01772_ _01773_ _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07098_ ci_neuron.uut_simple_neuron.x3\[22\] _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout232 net233 net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06049_ ci_neuron.uut_simple_neuron.x2\[27\] _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout221 net222 net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout210 net211 net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout243 net246 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07176__A1 _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout265 net266 net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout254 net258 net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout287 net288 net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout276 net283 net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09808_ _00387_ net42 internal_ih.byte7\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09739_ _00318_ net222 ci_neuron.uut_simple_neuron.x2\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08676__B2 _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09228__I0 _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout178_I net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05420_ _00969_ ci_neuron.uut_simple_neuron.x2\[13\] ci_neuron.uut_simple_neuron.x2\[14\]
+ _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_56_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05351_ _00999_ _01023_ _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_126_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05282_ _00954_ _00956_ _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_71_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08070_ _03621_ _03622_ _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09219__I0 _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07021_ _02599_ _02605_ _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08972_ internal_ih.byte7\[3\] internal_ih.byte6\[3\] _04332_ _04334_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07923_ ci_neuron.uut_simple_neuron.titan_id_2\[16\] ci_neuron.uut_simple_neuron.titan_id_5\[16\]
+ _03500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07854_ _03434_ _03435_ _03440_ _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06805_ _02387_ _02389_ _02442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_07785_ _03385_ _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_97_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04997_ internal_ih.byte2\[6\] _00691_ _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06736_ _02085_ _02343_ _02373_ _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_79_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09524_ _04721_ _04733_ _04735_ _04736_ _00538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06667_ _02306_ _00234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09455_ _03795_ ci_neuron.input_memory\[1\]\[12\] _00971_ _02226_ _04667_ _04669_
+ _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_66_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05618_ _01260_ _01284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08406_ _03909_ _00189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06598_ _02235_ _02238_ _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09386_ _04603_ _04618_ _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05549_ _01183_ _01194_ _01216_ _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_74_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08337_ _03848_ _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_22_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09473__I3 _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08268_ ci_neuron.uut_simple_neuron.x0\[11\] ci_neuron.uut_simple_neuron.x0\[12\]
+ _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__08425__A4 _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07219_ _02792_ _02832_ _02849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09485__I _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10230_ _00157_ net192 ci_neuron.uut_simple_neuron.titan_id_6\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08199_ ci_neuron.uut_simple_neuron.x0\[3\] _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07397__A1 _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_5_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10161_ _00077_ net197 ci_neuron.uut_simple_neuron.titan_id_2\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10092_ _00189_ net74 ci_neuron.uut_simple_neuron.titan_id_0\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_128_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08821__A1 _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04920_ _00649_ _00005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07560__A1 _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04851_ internal_ih.byte4\[0\] internal_ih.byte3\[0\] _00601_ _00602_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06259__I _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07570_ _00162_ _03129_ _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06521_ _02119_ _02163_ _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09240_ _04523_ _00467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06452_ _02001_ _02095_ _02096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_91_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07863__A2 ci_neuron.uut_simple_neuron.titan_id_5\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06383_ _02018_ _02019_ _02028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05403_ _01032_ _01063_ _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09171_ ci_neuron.uut_simple_neuron.titan_id_6\[29\] _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05334_ _00970_ _01006_ _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08812__A1 _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09455__I3 _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08122_ ci_neuron.uut_simple_neuron.titan_id_1\[19\] ci_neuron.uut_simple_neuron.titan_id_0\[19\]
+ _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_60_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08053_ _03608_ _00092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07004_ _02515_ _02517_ _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05265_ _00939_ _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05196_ _00855_ _00873_ _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08955_ _04324_ _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07906_ _03486_ _00131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08886_ _04269_ _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07837_ ci_neuron.uut_simple_neuron.titan_id_2\[2\] ci_neuron.uut_simple_neuron.titan_id_5\[2\]
+ _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07768_ _03368_ _03369_ _03371_ _03372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_27_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06719_ _02308_ _02357_ _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09507_ _04674_ _04722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_123_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07699_ ci_neuron.uut_simple_neuron.titan_id_4\[9\] ci_neuron.uut_simple_neuron.titan_id_3\[9\]
+ _03312_ _03313_ _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09438_ _04652_ _04662_ _04663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09369_ _03930_ _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08803__A1 _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09446__I3 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05093__A2 _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10213_ _00110_ net247 ci_neuron.uut_simple_neuron.titan_id_5\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_101_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10144_ _00209_ net286 ci_neuron.uut_simple_neuron.titan_id_3\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10075_ _00172_ net181 ci_neuron.uut_simple_neuron.titan_id_0\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08893__I1 internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07845__A2 ci_neuron.uut_simple_neuron.titan_id_5\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09437__I3 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08645__I1 ci_neuron.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06820__A3 _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05050_ _00734_ _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05952_ _00748_ _01582_ _01581_ _01610_ _01529_ _01611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_08740_ internal_ih.received_byte_count\[3\] _04197_ _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05883_ _01518_ _01520_ _01543_ _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XPHY_EDGE_ROW_77_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09373__I2 _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04903_ _00638_ _00022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08671_ spi_interface_cvonk.state\[1\] spi_interface_cvonk.state\[0\] _04139_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09522__A2 _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07622_ _00163_ _03206_ _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04834_ internal_ih.received_byte_count\[4\] internal_ih.received_byte_count\[7\]
+ internal_ih.received_byte_count\[6\] _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_109_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07553_ _02550_ _03178_ _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09286__A1 _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07484_ _02444_ _03025_ _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06504_ _02138_ _02146_ _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_76_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08884__I1 internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06435_ _01868_ _01954_ _02078_ _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__05847__A1 _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09223_ _04499_ _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_118_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_86_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09154_ _04473_ _00431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06366_ _01987_ _01993_ _02011_ _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_08105_ _03648_ _03649_ _03651_ _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_8_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08932__I _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06297_ _01909_ _01911_ _01944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05317_ _00960_ _00990_ _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09085_ _04415_ _04426_ _04428_ _00407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05248_ _00889_ _00899_ _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08036_ ci_neuron.uut_simple_neuron.titan_id_1\[6\] ci_neuron.uut_simple_neuron.titan_id_0\[6\]
+ _03594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05179_ _00835_ _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09987_ _00502_ net173 ci_neuron.input_memory\[1\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_95_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08938_ internal_ih.byte5\[4\] internal_ih.byte4\[4\] _04312_ _04315_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_4_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08869_ internal_ih.byte1\[6\] internal_ih.byte0\[6\] _04275_ _04276_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_125_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09277__A1 _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08875__I1 internal_ih.byte1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10127_ _00159_ net264 ci_neuron.uut_simple_neuron.titan_id_3\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10058_ _00543_ net137 ci_neuron.output_val_internal\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout258_I net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05829__A1 _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08866__I1 internal_ih.byte0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06220_ _01867_ _01861_ _01869_ _01870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08491__A2 _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06151_ _01785_ _01788_ _01805_ _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_13_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06272__I _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06082_ _01694_ _01722_ _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05102_ _00734_ _00770_ _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05033_ ci_neuron.address_i\[5\] ci_neuron.address_i\[4\] ci_neuron.address_i\[3\]
+ _00719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09910_ _00006_ net8 ci_neuron.address_i\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09841_ _00420_ net160 ci_neuron.output_memory\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06984_ _02615_ _02617_ _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_95_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09772_ _00351_ net49 internal_ih.byte2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout73_I net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05935_ _01515_ _01544_ _01595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08723_ _04179_ _04182_ _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05866_ _01526_ _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08654_ _04123_ _00281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05797_ _01437_ _01439_ _01459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07605_ ci_neuron.uut_simple_neuron.x3\[28\] _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08585_ _03838_ _04049_ _04066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_37_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07536_ _03160_ _03161_ _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_120_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07467_ _02727_ _02867_ _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09206_ _03770_ _04500_ _04505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07398_ _02444_ _03025_ _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06418_ _02062_ _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08609__I1 _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06349_ _01966_ _01995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09137_ ci_neuron.uut_simple_neuron.titan_id_6\[12\] _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09431__A1 ci_neuron.output_memory\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06245__A1 _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09068_ ci_neuron.stream_o\[27\] _04381_ _04412_ _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08019_ ci_neuron.uut_simple_neuron.titan_id_1\[2\] ci_neuron.uut_simple_neuron.titan_id_0\[2\]
+ _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08793__I0 _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05220__A2 _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08837__I _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05261__I _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09489__A1 ci_neuron.output_memory\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05720_ _01329_ _01380_ _01383_ _01384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05651_ _01283_ _01298_ _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_106_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08370_ _03877_ _03875_ _03878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07321_ _02924_ _02949_ _02950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_92_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05582_ _01217_ _01231_ _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08839__I1 _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08464__A2 _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07252_ _02341_ _02881_ _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07183_ _02494_ _02813_ _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06203_ _01853_ _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07098__I ci_neuron.uut_simple_neuron.x3\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06134_ _01762_ _01789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_112_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06065_ _01699_ _01721_ _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05016_ _00704_ _00056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09824_ _00403_ net131 internal_ih.spi_tx_byte_o\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06967_ _02131_ _02543_ _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09755_ _00334_ net124 internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06898_ _02047_ _02490_ _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05918_ _01472_ _01577_ _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09686_ _00273_ net92 ci_neuron.uut_simple_neuron.x3\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08706_ internal_ih.spi_rx_byte_i\[7\] _04166_ _04142_ _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05849_ _01510_ _00215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_68_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08637_ _04107_ _04108_ _04109_ _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_77_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout10 net12 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout21 net22 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08568_ _04048_ _04050_ _04051_ _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07519_ _03143_ _03144_ _03145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout54 net55 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout43 net52 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout32 net34 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout65 net71 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08455__A2 _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08499_ _03769_ _03987_ _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xfanout87 net88 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout98 net101 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout76 net78 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08766__I0 _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05432__A2 _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07870_ _03435_ _03440_ _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06821_ _02434_ _02457_ _02458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06752_ _02387_ _02389_ _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09540_ _04743_ _04745_ _04748_ _04750_ _00540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_92_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05703_ _00750_ _01329_ _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09471_ _04666_ _04691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06683_ _02045_ _02181_ _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08422_ ci_neuron.instruction_i\[2\] _03922_ _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_47_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05634_ _01067_ _01299_ _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05115__B _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05565_ _01215_ _01232_ _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08353_ ci_neuron.uut_simple_neuron.x0\[23\] _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07304_ _02734_ _02735_ _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06448__A1 _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08284_ ci_neuron.uut_simple_neuron.x0\[13\] ci_neuron.uut_simple_neuron.x0\[14\]
+ _03803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_05496_ _01075_ _01157_ _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07235_ ci_neuron.uut_simple_neuron.x3\[24\] _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_34_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07166_ ci_neuron.uut_simple_neuron.x3\[23\] _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07097_ _02548_ _02683_ _02728_ _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06117_ _01699_ _01721_ _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06048_ _01663_ _01703_ _01704_ _01621_ _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_100_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout222 net224 net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout211 net212 net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout200 net203 net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout244 net246 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07176__A2 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout233 net234 net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout255 net257 net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout288 net289 net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout277 net282 net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout266 net272 net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09807_ _00386_ net41 internal_ih.byte7\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07999_ _03541_ _03542_ _03559_ _03564_ _03565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_09738_ _00317_ net222 ci_neuron.uut_simple_neuron.x2\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ _00256_ net259 ci_neuron.uut_simple_neuron.x3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07939__A1 _03512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08987__I0 _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08600__A2 _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06678__A1 _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout240_I net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_44_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05350_ _01001_ _01004_ _01022_ _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_83_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05281_ _00927_ _00926_ _00928_ _00955_ _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_71_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07020_ _02602_ _02604_ _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08971_ _04333_ _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07922_ _03499_ _00134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07158__A2 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07853_ _03441_ _00154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06804_ _02386_ _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07784_ ci_neuron.uut_simple_neuron.titan_id_4\[24\] ci_neuron.uut_simple_neuron.titan_id_3\[24\]
+ ci_neuron.uut_simple_neuron.titan_id_4\[23\] ci_neuron.uut_simple_neuron.titan_id_3\[23\]
+ _03385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_97_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_04996_ _00693_ _00046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06735_ _02086_ _02222_ _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_79_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09523_ ci_neuron.output_val_internal\[22\] _04727_ _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06666_ _02303_ _02305_ _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_65_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09454_ _04602_ _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05617_ _01257_ _01274_ _01282_ _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09385_ _03724_ ci_neuron.input_memory\[1\]\[2\] _00774_ _01849_ _04605_ _04607_
+ _04618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08405_ _03904_ _03905_ _03908_ _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06597_ _02237_ _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_52_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08336_ ci_neuron.uut_simple_neuron.x0\[20\] _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05548_ _00751_ _01152_ _01193_ _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_62_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05479_ ci_neuron.uut_simple_neuron.x2\[16\] _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08267_ _03788_ _00171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07218_ _02792_ _02832_ _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06841__A1 _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08198_ _03728_ _00190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_120_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07149_ _02710_ _02711_ _02715_ _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07286__I _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09630__I1 ci_neuron.output_memory\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08594__A1 _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10160_ _00066_ net187 ci_neuron.uut_simple_neuron.titan_id_2\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10091_ _00188_ net76 ci_neuron.uut_simple_neuron.titan_id_0\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__04907__A1 internal_ih.byte5\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04907__B2 internal_ih.byte1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_106_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_127_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08821__A2 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_115_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10289_ _00582_ net139 ci_neuron.stream_o\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout288_I net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04850_ _00600_ _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05571__A1 _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_124_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06520_ _02120_ _02162_ _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08755__I _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06451_ _02090_ _02094_ _02095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05402_ _01073_ _00205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05323__A1 _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06382_ _01981_ _02023_ _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09170_ _04481_ _00439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05333_ _01005_ _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_60_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08121_ _03658_ _03663_ _03665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05264_ ci_neuron.uut_simple_neuron.x2\[9\] ci_neuron.uut_simple_neuron.x2\[10\]
+ ci_neuron.uut_simple_neuron.x2\[11\] _00939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_08052_ _03606_ _03607_ _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07003_ _02634_ _02636_ _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_113_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05195_ _00856_ _00872_ _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08954_ internal_ih.byte6\[3\] internal_ih.byte5\[3\] _04322_ _04324_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07905_ ci_neuron.uut_simple_neuron.titan_id_2\[13\] ci_neuron.uut_simple_neuron.titan_id_5\[13\]
+ _03485_ _03486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08885_ _04284_ _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07836_ ci_neuron.uut_simple_neuron.titan_id_2\[2\] ci_neuron.uut_simple_neuron.titan_id_5\[2\]
+ _03427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07767_ ci_neuron.uut_simple_neuron.titan_id_4\[21\] ci_neuron.uut_simple_neuron.titan_id_3\[21\]
+ _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_04979_ _00683_ _00038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06718_ _02355_ _02356_ _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09506_ _04696_ _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07698_ _03314_ _00125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08500__A1 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06649_ _02282_ _02288_ _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09437_ _04005_ ci_neuron.input_memory\[1\]\[10\] _00911_ _02091_ _04644_ _04645_
+ _04662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_19_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09368_ _04602_ _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09299_ ci_neuron.input_memory\[1\]\[10\] _04556_ _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08319_ _03832_ _03830_ _03831_ _03834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_35_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08803__A2 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10212_ _00109_ net243 ci_neuron.uut_simple_neuron.titan_id_5\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_120_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10143_ _00208_ net286 ci_neuron.uut_simple_neuron.titan_id_3\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10074_ _00171_ net205 ci_neuron.uut_simple_neuron.titan_id_0\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_54_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06805__A1 _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08524__B _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05951_ _01584_ _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05882_ _01538_ _01542_ _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_84_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09373__I3 _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04902_ internal_ih.byte4\[7\] _00633_ _00634_ internal_ih.byte0\[7\] _00638_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08670_ spi_interface_cvonk.SCLK_r\[2\] _04125_ _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07621_ _03203_ _03205_ _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04833_ _00583_ internal_ih.received_byte_count\[2\] internal_ih.expected_byte_count\[3\]
+ _00584_ _00585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07552_ _02559_ _03177_ _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_109_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06503_ _02045_ _02145_ _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_76_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07483_ _02451_ _03024_ _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06434_ _02055_ _02056_ _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09222_ _04513_ _00459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06365_ _02006_ _02010_ _02011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09153_ ci_neuron.uut_simple_neuron.titan_id_6\[20\] _04473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05316_ _00879_ _00989_ _00990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08104_ ci_neuron.uut_simple_neuron.titan_id_1\[16\] ci_neuron.uut_simple_neuron.titan_id_0\[16\]
+ _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_32_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06296_ _01912_ _01914_ _01941_ _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09084_ internal_ih.spi_tx_byte_o\[4\] _04427_ _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10218__CLK net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05247_ _00889_ _00899_ _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08035_ _03590_ _03592_ _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05178_ _00820_ _00853_ _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_73_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_73_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09210__A2 _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09986_ _00501_ net94 ci_neuron.input_memory\[1\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08937_ _04314_ _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08868_ _04269_ _04275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_125_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07819_ ci_neuron.uut_simple_neuron.titan_id_4\[30\] ci_neuron.uut_simple_neuron.titan_id_3\[30\]
+ _03414_ _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08799_ _04052_ _01184_ _04231_ _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09521__I0 _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06263__A2 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10126_ net38 net264 ci_neuron.uut_simple_neuron.titan_id_3\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10057_ _00542_ net137 ci_neuron.output_val_internal\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08779__A1 _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06150_ _01791_ _01804_ _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06081_ _01736_ _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05101_ _00781_ _00761_ _00782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05032_ ci_neuron.address_i\[17\] ci_neuron.address_i\[16\] ci_neuron.address_i\[15\]
+ ci_neuron.address_i\[14\] _00718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_1_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09683__CLK net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09840_ _00419_ net192 ci_neuron.output_memory\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06983_ _02616_ _02556_ _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09771_ _00350_ net65 internal_ih.byte2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05934_ _01236_ _01594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08722_ _04173_ _04174_ _04181_ _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_96_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05865_ _01374_ _01461_ _01525_ _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08653_ _04122_ ci_neuron.uut_simple_neuron.x3\[31\] _04111_ _04123_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05796_ _01426_ _01457_ _01458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07604_ _03084_ _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08584_ _04065_ _00269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07535_ _03093_ _03097_ _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_120_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07466_ _03082_ _03092_ _03093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06417_ _01985_ _02036_ _02061_ _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_107_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09205_ _03990_ _04503_ _04504_ _00451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04879__I0 internal_ih.byte4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07397_ _02451_ _03024_ _03025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06348_ _01963_ _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09136_ _04464_ _00422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06279_ _01925_ _01926_ _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09067_ _04382_ _04408_ _04410_ _04411_ _04412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_32_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08018_ _03579_ _00127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09969_ _00484_ net178 ci_neuron.input_memory\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05028__B _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07984__A2 ci_neuron.uut_simple_neuron.titan_id_5\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09186__A1 _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10109_ _00233_ net281 ci_neuron.uut_simple_neuron.titan_id_4\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05650_ _01315_ _00211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_106_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05581_ _01075_ _01234_ _01247_ _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_34_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07320_ _02945_ _02948_ _02949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08763__I _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07251_ _02494_ _02813_ _02880_ _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07182_ _02449_ _02812_ _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06202_ _01844_ _01853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06133_ _01786_ _01787_ _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08472__I0 _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07975__A2 ci_neuron.uut_simple_neuron.titan_id_5\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06064_ _01702_ _01720_ _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_41_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05015_ internal_ih.byte3\[6\] _00701_ _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09823_ _00402_ net132 internal_ih.instruction_received vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06966_ _02132_ _02542_ _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09754_ _00333_ net60 internal_ih.byte0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06897_ _02082_ _02489_ _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09685_ _00272_ net226 ci_neuron.uut_simple_neuron.x3\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05917_ ci_neuron.uut_simple_neuron.x2\[25\] ci_neuron.uut_simple_neuron.x2\[26\]
+ _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_08705_ _04147_ _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05848_ _01495_ _01509_ _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08636_ ci_neuron.value_i\[28\] _04001_ _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05779_ _01415_ _01441_ _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_81_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout11 net12 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout22 net26 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08567_ ci_neuron.value_i\[17\] _04032_ _04051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07518_ _03066_ _03141_ _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08498_ _03986_ _03990_ _03991_ _00257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout55 net56 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout44 net46 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout33 net34 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07449_ _03004_ _03021_ _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_107_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout88 net91 net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout66 net71 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout77 net78 net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout99 net101 net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07415__A1 _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09119_ ci_neuron.uut_simple_neuron.titan_id_6\[3\] _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05977__A1 _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08766__I1 _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09009__I internal_ih.data_pointer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07654__A1 ci_neuron.uut_simple_neuron.titan_id_4\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07957__A2 ci_neuron.uut_simple_neuron.titan_id_5\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06820_ _02438_ _02440_ _02456_ _02457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__08758__I _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06751_ ci_neuron.uut_simple_neuron.x3\[16\] _02388_ _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_92_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06682_ _02275_ _02294_ _02320_ _02321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05702_ _01362_ _01364_ _01365_ _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_19_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09470_ ci_neuron.output_memory\[15\] _04675_ _04690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08421_ _00711_ _00712_ _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05633_ _01283_ _01298_ _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09589__I _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05564_ _01217_ _01231_ _01232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09871__CLK net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08352_ _03861_ _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07303_ _02727_ _02871_ _02931_ _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06448__A2 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05495_ _01126_ _01156_ _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08283_ _03802_ _00173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07234_ _02797_ _02863_ _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_63_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_119_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09398__A1 ci_neuron.output_memory\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07165_ _02739_ _02741_ _02795_ _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07096_ _02725_ _02727_ _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06116_ _01702_ _01720_ _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06047_ _01668_ _01622_ _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout223 net224 net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout212 net213 net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout201 net203 net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout245 net248 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout256 net257 net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout234 net252 net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout289 net290 net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout278 net282 net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout267 net271 net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09806_ _00385_ net42 internal_ih.byte6\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07998_ ci_neuron.uut_simple_neuron.titan_id_2\[27\] ci_neuron.uut_simple_neuron.titan_id_5\[27\]
+ _03558_ _03561_ _03563_ _03564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06949_ _02357_ _02410_ _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09737_ _00316_ net227 ci_neuron.uut_simple_neuron.x2\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09668_ _00255_ net259 ci_neuron.uut_simple_neuron.x3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08619_ _04094_ _02934_ _04086_ _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09599_ _04789_ _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_108_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06916__I ci_neuron.uut_simple_neuron.x3\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__A2 _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09389__A1 ci_neuron.output_memory\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout233_I net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05280_ _00922_ _00925_ _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06850__A2 _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08970_ internal_ih.byte7\[2\] internal_ih.byte6\[2\] _04332_ _04333_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07921_ _03497_ _03498_ _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07852_ _03439_ _03440_ _03441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06803_ _02393_ _02396_ _02439_ _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xinput1 spi_clock_i net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07783_ _03377_ _03382_ _03384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04995_ internal_ih.byte2\[5\] _00691_ _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09522_ _04724_ _04734_ _04735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06734_ _02325_ _02370_ _02371_ _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06665_ _02250_ _02253_ _02304_ _02305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09453_ ci_neuron.output_memory\[12\] _04675_ _04676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05616_ _01259_ _01273_ _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09384_ ci_neuron.output_memory\[2\] _04600_ _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08404_ _03906_ _03907_ _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06596_ _01994_ _02236_ _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08335_ _03847_ _00180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05547_ _01105_ _01209_ _01182_ _01214_ _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_47_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05478_ _01097_ _01147_ _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08266_ _03782_ _03785_ _03787_ _03788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_50_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06841__A2 _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07217_ _02787_ _02788_ _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08197_ _03724_ _03727_ _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07148_ _02761_ _02763_ _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07079_ _02661_ _02667_ _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10090_ _00187_ net77 ci_neuron.uut_simple_neuron.titan_id_0\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10124__CLK net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10288_ _00581_ net136 ci_neuron.stream_o\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09534__A1 ci_neuron.output_memory\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06450_ ci_neuron.uut_simple_neuron.x3\[11\] _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05401_ _01071_ _01072_ _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08972__S _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06381_ _01981_ _02023_ _02025_ _02026_ _00228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_84_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05332_ ci_neuron.uut_simple_neuron.x2\[13\] _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_60_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08120_ _03664_ _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05263_ _00937_ _00916_ _00938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08051_ ci_neuron.uut_simple_neuron.titan_id_1\[8\] ci_neuron.uut_simple_neuron.titan_id_0\[8\]
+ _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07002_ _02526_ _02568_ _02635_ _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_114_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05194_ _00841_ _00853_ _00871_ _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_12_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08953_ _04323_ _00380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07904_ _03481_ _03482_ _03484_ _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09525__A1 ci_neuron.output_memory\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06339__A1 _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08884_ internal_ih.byte2\[5\] internal_ih.byte1\[5\] _04280_ _04284_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05011__A1 internal_ih.byte3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07835_ _03426_ _00149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07766_ _03370_ _00108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04978_ internal_ih.byte1\[6\] _00680_ _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06717_ _02257_ _02299_ _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_79_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09505_ _04697_ _04715_ _04719_ _04720_ _00535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_93_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07697_ _03312_ _03313_ _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09436_ ci_neuron.output_memory\[10\] _04650_ _04661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06648_ _02144_ _02287_ _02288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_93_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06579_ _02184_ _02190_ _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08639__I0 _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09367_ _00728_ _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09298_ _04559_ _00489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08318_ _03830_ _03831_ _03832_ _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08249_ _03756_ _03769_ _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10211_ _00108_ net243 ci_neuron.uut_simple_neuron.titan_id_5\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10142_ _00207_ net286 ci_neuron.uut_simple_neuron.titan_id_3\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10073_ _00170_ net203 ci_neuron.uut_simple_neuron.titan_id_0\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05002__A1 internal_ih.byte3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07935__I _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05950_ _01526_ _01586_ _01608_ _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05881_ _01252_ _01254_ _01541_ _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_04901_ _00637_ _00021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07620_ _03243_ _03244_ _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04832_ internal_ih.received_byte_count\[3\] _00584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07551_ _02725_ _03096_ _03095_ _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_109_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06502_ _02141_ _02144_ _02145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_88_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08869__I0 internal_ih.byte1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07482_ _03107_ _03108_ _03109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_122_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06433_ _02039_ _02060_ _02076_ _02077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09221_ _04040_ _03825_ _04509_ _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06364_ _02009_ _02010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09152_ _04472_ _00430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05315_ _00946_ _00988_ _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08103_ _03650_ _00071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06295_ _01942_ _00168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09083_ _04377_ _04427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05246_ _00905_ _00921_ _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08034_ _03588_ _03591_ _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05177_ _00735_ _00838_ _00833_ _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_73_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09597__I1 ci_neuron.output_memory\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09985_ _00500_ net93 ci_neuron.input_memory\[1\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08936_ internal_ih.byte5\[3\] internal_ih.byte4\[3\] _04312_ _04314_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08867_ _04274_ _00343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07818_ _03410_ _03412_ _03413_ _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06732__A1 _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08798_ _04234_ _00314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07749_ _03348_ _03353_ _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07288__A2 _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08485__A1 _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09521__I1 ci_neuron.input_memory\[1\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09419_ _04630_ _04646_ _04647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_81_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07755__I _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10125_ _00249_ net235 ci_neuron.uut_simple_neuron.titan_id_4\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10056_ _00541_ net136 ci_neuron.output_val_internal\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08712__A2 _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08476__A1 ci_neuron.value_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06080_ _01734_ _01735_ _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05100_ net38 _00781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_13_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05031_ ci_neuron.address_i\[13\] ci_neuron.address_i\[12\] ci_neuron.address_i\[11\]
+ ci_neuron.address_i\[10\] _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_95_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07754__A3 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06982_ _02498_ _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09770_ _00349_ net63 internal_ih.byte2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05933_ _01449_ _01592_ _01593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08721_ internal_ih.instruction_received internal_ih.spi_rx_byte_i\[3\] _04180_ _04181_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_28_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08652_ ci_neuron.value_i\[31\] _04121_ _04026_ _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07603_ _03226_ _03227_ _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05864_ _01327_ _01524_ _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_89_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05795_ _01432_ _01436_ _01457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08583_ _04064_ _02552_ _04053_ _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07534_ _03082_ _03092_ _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07465_ _02870_ _03091_ _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_119_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06416_ _02039_ _02060_ _02061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09204_ _03756_ _04500_ _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07396_ _02615_ _03022_ _03023_ _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06347_ _01989_ _01990_ _01992_ _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09135_ ci_neuron.uut_simple_neuron.titan_id_6\[11\] _04464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06278_ _01905_ _01926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09066_ _04182_ _04411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05229_ _00787_ _00836_ _00904_ _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08017_ ci_neuron.uut_simple_neuron.titan_id_2\[0\] ci_neuron.uut_simple_neuron.titan_id_5\[0\]
+ _03579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09968_ _00483_ net178 ci_neuron.input_memory\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09578__S0 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08919_ internal_ih.byte4\[4\] internal_ih.byte3\[4\] _04301_ _04304_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09899_ _00018_ net10 ci_neuron.address_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09498__A3 _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05444__A1 _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07197__A1 _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09186__A2 _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10108_ _00232_ net281 ci_neuron.uut_simple_neuron.titan_id_4\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10039_ _00524_ net169 ci_neuron.output_val_internal\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout263_I net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05580_ _01206_ _01233_ _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08449__A1 _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07250_ _02495_ _02812_ _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08980__S _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07181_ _02622_ _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06201_ _01842_ _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07424__A2 _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06132_ _01450_ _01777_ _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08472__I1 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06063_ _01661_ _01719_ _01720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05014_ _00703_ _00054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09822_ _00401_ net57 internal_ih.current_instruction\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09753_ _00332_ net122 internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06965_ _02597_ _02598_ _02599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08704_ _04133_ _04164_ _04165_ _00289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06896_ _02529_ _02530_ _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05916_ _00937_ _01575_ _01569_ _01576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09684_ _00271_ net226 ci_neuron.uut_simple_neuron.x3\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05847_ _01500_ _01502_ _01508_ _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_49_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08635_ _03904_ _04106_ _03959_ _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_68_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08566_ _03971_ _04049_ _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07517_ _03068_ _03140_ _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05778_ _01418_ _01440_ _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_81_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout12 net17 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08497_ _01961_ _03980_ _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout56 net62 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout34 net35 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout23 net25 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout45 net46 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07448_ _03028_ _03038_ _03074_ _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout89 net90 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout67 net70 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout78 net79 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07379_ _03005_ _03006_ _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09118_ _04455_ _00413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09049_ internal_ih.spi_tx_byte_o\[1\] _04379_ _04396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05665__A1 _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06750_ ci_neuron.uut_simple_neuron.x3\[17\] _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06681_ _02278_ _02293_ _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05701_ _01331_ _01363_ _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_19_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07342__A1 _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05632_ _01284_ _01297_ _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08420_ _03921_ _00192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_47_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05563_ _01221_ _01230_ _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08351_ ci_neuron.uut_simple_neuron.x0\[22\] _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07302_ _02930_ _02870_ _02931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05494_ _01163_ _00207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08282_ _03798_ _03801_ _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08842__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07233_ ci_neuron.uut_simple_neuron.x3\[24\] _02863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05656__A1 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07164_ _02729_ _02738_ _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_6_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07095_ _02726_ _02681_ _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06115_ _01698_ _01746_ _01770_ _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06046_ _01672_ _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout213 net214 net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout202 net203 net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout246 net248 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout235 net236 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout224 net225 net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout279 net281 net279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout257 net258 net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout268 net271 net268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09805_ _00384_ net40 internal_ih.byte6\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07997_ _03562_ _03563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06948_ _02578_ _02579_ _02580_ _02582_ _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_09736_ _00315_ net226 ci_neuron.uut_simple_neuron.x2\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09667_ _00254_ net259 ci_neuron.uut_simple_neuron.x3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06879_ _02472_ _02514_ _02515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08618_ _04091_ _04093_ _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09720__D _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09598_ _04794_ _00554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08549_ _04035_ _00264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__C _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07636__A2 _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08859__I _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09400__I3 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04861__A2 _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07920_ ci_neuron.uut_simple_neuron.titan_id_2\[16\] ci_neuron.uut_simple_neuron.titan_id_5\[16\]
+ _03498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07851_ ci_neuron.uut_simple_neuron.titan_id_2\[5\] ci_neuron.uut_simple_neuron.titan_id_5\[5\]
+ _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06802_ _02382_ _02392_ _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07782_ _03383_ _00111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06366__A2 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput2 spi_cs_i net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06733_ _02328_ _02346_ _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09521_ _03862_ ci_neuron.input_memory\[1\]\[22\] _01381_ _02805_ _04716_ _04717_
+ _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_04994_ _00692_ _00045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06664_ _02209_ _02249_ _02304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_65_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09452_ _04674_ _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05615_ _01281_ _00210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06595_ _01995_ _02093_ _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_09383_ _04598_ _04613_ _04615_ _04616_ _00517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_08403_ _03898_ _03901_ _03907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05546_ _01212_ _01213_ _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08334_ _03844_ _03846_ _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_22_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05477_ _01146_ _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08265_ _03777_ _03780_ _03786_ _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07216_ _02835_ _02838_ _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08196_ _03725_ _03726_ _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07147_ _02774_ _02776_ _02777_ _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_104_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06054__A1 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07078_ _02664_ _02666_ _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06029_ _01686_ _00219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09543__A2 _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09719_ _00298_ net255 ci_neuron.uut_simple_neuron.x2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10287_ _00580_ net140 ci_neuron.stream_o\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09385__I2 _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_49_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout176_I net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07442__B _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07848__A2 ci_neuron.uut_simple_neuron.titan_id_5\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05400_ _01029_ _01027_ _01070_ _01072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_56_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_38_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06380_ _02024_ _02023_ _02026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_83_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05331_ _00743_ _01002_ _00974_ _01003_ _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_60_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09470__A1 ci_neuron.output_memory\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05262_ _00936_ _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08050_ _03602_ _03603_ _03604_ _03605_ _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_3_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07001_ _02528_ _02567_ _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05193_ _00862_ _00870_ _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08952_ internal_ih.byte6\[2\] internal_ih.byte5\[2\] _04322_ _04323_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_47_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07903_ ci_neuron.uut_simple_neuron.titan_id_2\[12\] ci_neuron.uut_simple_neuron.titan_id_5\[12\]
+ _03484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08883_ _04283_ _00350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_71_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07834_ ci_neuron.uut_simple_neuron.titan_id_2\[2\] ci_neuron.uut_simple_neuron.titan_id_5\[2\]
+ _03425_ _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_127_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07765_ _03368_ _03369_ _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09289__A1 _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04977_ _00682_ _00037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06716_ _02309_ _02354_ _02355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07696_ ci_neuron.uut_simple_neuron.titan_id_4\[9\] ci_neuron.uut_simple_neuron.titan_id_3\[9\]
+ _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09504_ ci_neuron.output_val_internal\[19\] _04705_ _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06647_ _02285_ _02286_ _02287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_78_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_56_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08887__I1 internal_ih.byte1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09435_ _04649_ _04657_ _04659_ _04660_ _00525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_109_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06578_ _01870_ _02218_ _02219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09366_ ci_neuron.output_memory\[0\] _04600_ _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05529_ _01169_ _01197_ _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09297_ _04003_ ci_neuron.input_memory\[1\]\[9\] _04543_ _04559_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08317_ ci_neuron.uut_simple_neuron.x0\[17\] ci_neuron.uut_simple_neuron.x0\[18\]
+ _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_35_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08248_ _03771_ _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10210_ _00106_ net244 ci_neuron.uut_simple_neuron.titan_id_5\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_08179_ ci_neuron.uut_simple_neuron.titan_id_1\[29\] ci_neuron.uut_simple_neuron.titan_id_0\[29\]
+ _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_65_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10141_ _00206_ net280 ci_neuron.uut_simple_neuron.titan_id_3\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10072_ _00199_ net204 ci_neuron.uut_simple_neuron.titan_id_0\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08878__I1 internal_ih.byte1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04900_ internal_ih.byte4\[6\] _00633_ _00634_ internal_ih.byte0\[6\] _00637_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05880_ _01429_ _01539_ _01540_ _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_04831_ internal_ih.expected_byte_count\[2\] _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07550_ _03175_ _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_109_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06501_ _02090_ _02143_ _02144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08869__I1 internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07481_ _02041_ _03035_ _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09220_ _04512_ _00458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_122_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06432_ _02043_ _02059_ _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06363_ _02008_ _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09151_ ci_neuron.uut_simple_neuron.titan_id_6\[19\] _04472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05314_ _00962_ _00987_ _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08102_ _03648_ _03649_ _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09082_ ci_neuron.stream_o\[28\] _04416_ _04425_ _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_32_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06294_ _01916_ _01941_ _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08033_ ci_neuron.uut_simple_neuron.titan_id_1\[5\] ci_neuron.uut_simple_neuron.titan_id_0\[5\]
+ _03591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_4_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05245_ _00907_ _00920_ _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05176_ _00798_ _00818_ _00853_ _00843_ _00834_ _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_73_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09984_ _00499_ net93 ci_neuron.input_memory\[1\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10114__CLK net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08935_ _04313_ _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08866_ internal_ih.byte1\[5\] internal_ih.byte0\[5\] _04270_ _04274_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07817_ ci_neuron.uut_simple_neuron.titan_id_4\[29\] ci_neuron.uut_simple_neuron.titan_id_3\[29\]
+ _03413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_98_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08797_ _04046_ _01150_ _04231_ _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07748_ ci_neuron.uut_simple_neuron.titan_id_4\[18\] ci_neuron.uut_simple_neuron.titan_id_3\[18\]
+ _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_94_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07679_ ci_neuron.uut_simple_neuron.titan_id_4\[6\] ci_neuron.uut_simple_neuron.titan_id_3\[6\]
+ ci_neuron.uut_simple_neuron.titan_id_4\[5\] ci_neuron.uut_simple_neuron.titan_id_3\[5\]
+ _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__09521__I2 _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09418_ _03756_ ci_neuron.input_memory\[1\]\[7\] _00847_ _01961_ _04644_ _04645_
+ _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_51_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09349_ _04375_ internal_ih.expected_byte_count\[0\] _04353_ _04588_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_73_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05471__A2 _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10124_ _00248_ net241 ci_neuron.uut_simple_neuron.titan_id_4\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06971__A2 _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08548__I0 _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10055_ _00540_ net165 ci_neuron.output_val_internal\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_82_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06487__A1 _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_91_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05030_ ci_neuron.address_i\[21\] ci_neuron.address_i\[20\] ci_neuron.address_i\[19\]
+ ci_neuron.address_i\[18\] _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__08978__S _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06981_ _02554_ _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08539__I0 ci_neuron.value_i\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05932_ _01556_ _01591_ _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08720_ _04171_ _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05863_ _01342_ ci_neuron.uut_simple_neuron.x2\[22\] ci_neuron.uut_simple_neuron.x2\[23\]
+ _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08651_ ci_neuron.uut_simple_neuron.x0\[31\] _03920_ _04114_ _04121_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07602_ _03172_ _03173_ _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05794_ _01413_ _01454_ _01455_ _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08582_ _04061_ _04062_ _04063_ _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_37_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07533_ _03100_ _03103_ _03158_ _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07464_ _03090_ _03091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08726__B _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06415_ _02043_ _02059_ _02060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_57_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09203_ _04488_ _04503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07395_ _02557_ _02808_ _03023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09134_ _04463_ _00421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06346_ _01991_ _01969_ _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06277_ _01902_ _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09065_ _04389_ _04409_ _04410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05228_ _00833_ _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08016_ _03578_ _00151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08461__B _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05159_ _00837_ _00838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09967_ _00482_ net180 ci_neuron.input_memory\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09578__S1 _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08918_ _04303_ _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09898_ _00017_ net15 ci_neuron.address_i\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08849_ _04257_ _04264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_95_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09311__I _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05141__A1 _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10107_ _00231_ net286 ci_neuron.uut_simple_neuron.titan_id_4\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10038_ _00523_ net171 ci_neuron.output_val_internal\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08449__A2 _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06200_ _01836_ _01839_ _01851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_14_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07180_ _02803_ _02810_ _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_109_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06131_ _01740_ _01776_ _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06062_ _01705_ _01718_ _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_57_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05013_ internal_ih.byte3\[5\] _00701_ _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09821_ _00400_ net57 internal_ih.current_instruction\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09752_ _00331_ net60 internal_ih.byte0\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06964_ _01833_ _02535_ _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08703_ internal_ih.spi_rx_byte_i\[7\] _04148_ _04165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06895_ _01824_ _02481_ _02530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09683_ _00270_ net250 ci_neuron.uut_simple_neuron.x3\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05915_ _01574_ _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05846_ _01445_ _01504_ _01506_ _01507_ _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08634_ _03903_ _04106_ _04107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_05777_ _01437_ _01439_ _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_68_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08565_ _03824_ _04043_ _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07516_ _03142_ _00247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout13 net16 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout35 net36 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout24 net26 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout46 net47 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08496_ ci_neuron.value_i\[7\] _03952_ _03989_ _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_07447_ _03001_ _03027_ _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout57 net59 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout68 net70 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout79 net84 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07378_ _02863_ _02938_ _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06329_ _01945_ _01972_ _01975_ _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_60_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09117_ ci_neuron.uut_simple_neuron.titan_id_6\[2\] _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06623__A1 _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09048_ ci_neuron.stream_o\[25\] _04381_ _04394_ _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05362__A1 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07103__A2 ci_neuron.uut_simple_neuron.x3\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06680_ _02315_ _02318_ _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05700_ _01331_ _01363_ _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05631_ _01286_ _01296_ _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08350_ _03860_ _00182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_47_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07301_ _02927_ _02800_ _02929_ _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05562_ _01222_ _01229_ _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_74_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05493_ _01123_ _01162_ _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08281_ _03785_ _03799_ _03800_ _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08842__A2 _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07232_ _02625_ _02860_ _02861_ _02862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07163_ _02743_ _02747_ _02793_ _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_82_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06114_ _01700_ _01769_ _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_41_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07094_ _02620_ _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06045_ _01665_ _01673_ _01701_ _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05959__A3 _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout214 net215 net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout203 net207 net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08358__A1 _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout247 net249 net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout236 net242 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07030__A1 _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06908__A2 _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout225 net234 net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09804_ _00383_ net39 internal_ih.byte6\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout269 net271 net269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout258 net263 net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__04919__B2 internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07996_ ci_neuron.uut_simple_neuron.titan_id_2\[27\] ci_neuron.uut_simple_neuron.titan_id_5\[27\]
+ ci_neuron.uut_simple_neuron.titan_id_2\[26\] ci_neuron.uut_simple_neuron.titan_id_5\[26\]
+ _03562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06947_ _02521_ _02581_ _02582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09735_ _00314_ net228 ci_neuron.uut_simple_neuron.x2\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09666_ _00253_ net259 ci_neuron.uut_simple_neuron.x3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06878_ _02474_ _02513_ _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08617_ _03893_ _04082_ _04092_ _03959_ _04093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_05829_ _01078_ _01490_ _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09597_ ci_neuron.stream_o\[3\] ci_neuron.output_memory\[3\] _04790_ _04794_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08548_ _04034_ _02335_ _04028_ _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08479_ _03957_ _03974_ _03975_ _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08597__A1 _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08521__A1 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09321__I0 _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08824__A2 _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08588__A1 _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09624__I1 ci_neuron.output_memory\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07850_ _03437_ _03438_ _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07781_ _03381_ _03382_ _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06801_ _02040_ _02437_ _02438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08760__A1 _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04993_ internal_ih.byte2\[4\] _00691_ _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06732_ _02328_ _02346_ _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput3 spi_pico_i net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09520_ ci_neuron.output_memory\[22\] _04722_ _04733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06663_ _02301_ _02302_ _02303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09451_ _00727_ _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06594_ _02225_ _02234_ _02235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05614_ _01278_ _01280_ _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_93_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout34_I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09382_ ci_neuron.output_val_internal\[1\] _04611_ _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08402_ _03891_ _03903_ _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07079__A1 _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05545_ _00888_ _01142_ _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09312__I0 _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08333_ _03823_ _03835_ _03833_ _03837_ _03845_ _03846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_117_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08264_ _03771_ ci_neuron.uut_simple_neuron.x0\[10\] _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05476_ _01145_ _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07215_ _02843_ _02844_ _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09615__I1 ci_neuron.output_memory\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08195_ _00706_ _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07146_ _02583_ _02775_ _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07077_ _02656_ _02696_ _02708_ _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_76_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06028_ _01647_ _01685_ _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09718_ _00297_ net148 internal_ih.received_byte_count\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07979_ _03541_ _03542_ _03547_ _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07306__A2 _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08503__A1 _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09649_ _04823_ _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06293__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09606__I1 ci_neuron.output_memory\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08990__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04851__I0 internal_ih.byte4\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10286_ _00579_ net136 ci_neuron.stream_o\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09385__I3 _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_29_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05330_ _00968_ _00985_ _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07481__A1 _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05261_ _00747_ _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07000_ _02593_ _02596_ _02633_ _02634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_98_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05192_ _00835_ _00864_ _00869_ _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_102_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08951_ _04311_ _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07902_ _03483_ _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08882_ internal_ih.byte2\[4\] internal_ih.byte1\[4\] _04280_ _04283_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_71_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07833_ _03421_ _03422_ _03424_ _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_127_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07764_ ci_neuron.uut_simple_neuron.titan_id_4\[21\] ci_neuron.uut_simple_neuron.titan_id_3\[21\]
+ _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04976_ internal_ih.byte1\[5\] _00680_ _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06715_ _02351_ _02353_ _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07695_ _03308_ _03309_ _03310_ _03311_ _03312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_09503_ _04701_ _04718_ _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06646_ _02227_ ci_neuron.uut_simple_neuron.x3\[14\] ci_neuron.uut_simple_neuron.x3\[15\]
+ _02286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_94_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09434_ ci_neuron.output_val_internal\[9\] _04655_ _04660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_111_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06577_ _01882_ _02217_ _02218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09365_ _04599_ _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05528_ _01170_ _01196_ _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09296_ _03994_ _04553_ _04558_ _00488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08316_ _03810_ _03823_ _03821_ _03831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__06275__A2 _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05459_ _00961_ _01127_ _01128_ _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08247_ ci_neuron.uut_simple_neuron.x0\[9\] _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08178_ _03705_ _03710_ _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09213__A2 _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07129_ _02707_ _02709_ _02760_ _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XPHY_EDGE_ROW_120_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10140_ _00205_ net279 ci_neuron.uut_simple_neuron.titan_id_3\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10071_ _00198_ net202 ci_neuron.uut_simple_neuron.titan_id_0\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10269_ _00562_ net152 ci_neuron.stream_o\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07480_ _02436_ _02454_ _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_109_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06500_ ci_neuron.uut_simple_neuron.x3\[11\] _02142_ _02143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_119_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06431_ _00162_ _02074_ _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06362_ _01852_ _02007_ _02008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09150_ _04471_ _00429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06293_ _01919_ _01940_ _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05313_ _00966_ _00986_ _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08101_ ci_neuron.uut_simple_neuron.titan_id_1\[16\] ci_neuron.uut_simple_neuron.titan_id_0\[16\]
+ _03649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09081_ _04382_ _04422_ _04424_ _04411_ _04425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_32_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05244_ _00908_ _00919_ _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08032_ ci_neuron.uut_simple_neuron.titan_id_1\[5\] ci_neuron.uut_simple_neuron.titan_id_0\[5\]
+ _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05175_ _00840_ _00841_ _00852_ _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_101_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09983_ _00498_ net109 ci_neuron.input_memory\[1\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08934_ internal_ih.byte5\[2\] internal_ih.byte4\[2\] _04312_ _04313_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_4_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08865_ _04273_ _00342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07816_ ci_neuron.uut_simple_neuron.titan_id_4\[29\] ci_neuron.uut_simple_neuron.titan_id_3\[29\]
+ _03412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_98_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08796_ _04233_ _00313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07747_ _03354_ _00104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04959_ _00672_ _00060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10220__D _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07678_ _03287_ _03296_ _03297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09521__I3 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06629_ _02221_ _02239_ _02269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09417_ _04606_ _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09348_ _04587_ _00511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_51_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09279_ _03955_ _04544_ _04548_ _00481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07996__A2 ci_neuron.uut_simple_neuron.titan_id_5\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10123_ _00247_ net235 ci_neuron.uut_simple_neuron.titan_id_4\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08548__I1 _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10054_ _00539_ net167 ci_neuron.output_val_internal\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09044__I internal_ih.data_pointer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07987__A2 ci_neuron.uut_simple_neuron.titan_id_5\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06980_ _02560_ _02563_ _02613_ _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_95_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05931_ _01560_ _01590_ _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05862_ _01521_ _01484_ _01522_ _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08650_ _04120_ _00280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07601_ _03165_ _03171_ _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05793_ _01412_ _01438_ _01455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08581_ ci_neuron.value_i\[19\] _04032_ _04063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07532_ _03080_ _03098_ _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07463_ _03087_ _03089_ _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_76_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06414_ _02054_ _02058_ _02059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09202_ _03984_ _04494_ _04502_ _00450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07394_ _02557_ _02808_ _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09133_ ci_neuron.uut_simple_neuron.titan_id_6\[10\] _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06345_ _01957_ _01991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06276_ _01921_ _01922_ _01923_ _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09064_ ci_neuron.output_val_internal\[27\] ci_neuron.output_val_internal\[19\] ci_neuron.output_val_internal\[11\]
+ ci_neuron.output_val_internal\[3\] _04390_ _04391_ _04409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07978__A2 ci_neuron.uut_simple_neuron.titan_id_5\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05227_ _00903_ _00227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08015_ ci_neuron.uut_simple_neuron.titan_id_2\[31\] ci_neuron.uut_simple_neuron.titan_id_5\[31\]
+ _03577_ _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_05158_ _00833_ _00836_ _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05089_ _00734_ _00765_ _00770_ _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09966_ _00481_ net200 ci_neuron.input_memory\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08917_ internal_ih.byte4\[3\] internal_ih.byte3\[3\] _04301_ _04303_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09897_ _00012_ net14 ci_neuron.address_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08848_ _04263_ _00335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08779_ _03994_ _04218_ _04223_ _00306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07969__A2 ci_neuron.uut_simple_neuron.titan_id_5\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10106_ _00230_ net279 ci_neuron.uut_simple_neuron.titan_id_4\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10037_ _00522_ net170 ci_neuron.output_val_internal\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_106_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout151_I net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout249_I net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06130_ _01783_ _01784_ _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06061_ _01663_ _01717_ _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05012_ _00702_ _00053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09820_ _00399_ net58 internal_ih.current_instruction\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09582__A1 _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06963_ _02121_ _02103_ _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09751_ _00330_ net57 internal_ih.byte0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05914_ _01475_ _01573_ _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08702_ internal_ih.spi_tx_byte_o\[6\] _04136_ _04157_ internal_ih.spi_rx_byte_i\[6\]
+ _04164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06894_ _02074_ _02480_ _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09682_ _00269_ net226 ci_neuron.uut_simple_neuron.x3\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05845_ _01408_ _01503_ _01507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08633_ _03900_ _04102_ _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05776_ _01389_ _01438_ _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05371__A2 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08564_ _03840_ _04044_ _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07515_ _03066_ _03141_ _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout36 internal_ih.got_all_data net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout14 net16 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout47 net51 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout25 net26 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08495_ _03951_ _03987_ _03988_ _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_07446_ _03040_ _03053_ _03072_ _03073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout58 net61 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout69 net70 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07377_ _02868_ _02937_ _03005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06328_ _01920_ _01973_ _01974_ _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_32_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09116_ _04454_ _00412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06623__A2 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09047_ _04382_ _04388_ _04393_ _04354_ _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06259_ _01907_ _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_92_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09949_ _00464_ net99 ci_neuron.uut_simple_neuron.x0\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05630_ _01261_ _01295_ _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09232__I _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07300_ _02928_ _02865_ _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05561_ _01225_ _01228_ _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06302__A1 _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05492_ _01158_ _01161_ _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08280_ _03789_ _03792_ _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07231_ _02858_ _02859_ _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_63_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07162_ _02724_ _02742_ _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06113_ _01749_ _01768_ _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07093_ _02680_ _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08850__I0 internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06044_ _01700_ _01675_ _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08512__S _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout204 net206 net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout237 net240 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout226 net227 net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout215 net216 net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09803_ _00382_ net53 internal_ih.byte6\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout248 net249 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout259 net262 net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07995_ _03547_ _03560_ _03545_ _03561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06946_ _02522_ _02581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09734_ _00313_ net230 ci_neuron.uut_simple_neuron.x2\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06877_ _02484_ _02512_ _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09665_ _00252_ net275 ci_neuron.uut_simple_neuron.x3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05828_ _01453_ _01489_ _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08616_ _03876_ _03879_ _04082_ _04092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09596_ _04793_ _00553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05759_ _01375_ _01337_ _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_65_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08547_ _03952_ _04031_ _04033_ _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_119_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08478_ _01874_ _03948_ _03975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07429_ _02920_ _02972_ _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09546__A1 ci_neuron.output_memory\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08521__A2 _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout114_I net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07780_ ci_neuron.uut_simple_neuron.titan_id_4\[24\] ci_neuron.uut_simple_neuron.titan_id_3\[24\]
+ _03382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06800_ _02005_ _02436_ _02437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04992_ _00685_ _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput4 sys_clock_i net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06731_ _02316_ _02368_ _02369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08899__I0 internal_ih.byte3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09450_ _04597_ _04673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06662_ _02244_ _02255_ _02300_ _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_65_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08401_ ci_neuron.uut_simple_neuron.x0\[29\] _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06593_ _02136_ _02233_ _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05613_ _01240_ _01245_ _01279_ _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09381_ _04603_ _04614_ _04615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05544_ _01210_ _01211_ _01212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08332_ _03838_ _03845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout27_I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08263_ _03784_ _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07214_ _02778_ _02841_ _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05475_ _01099_ _01102_ _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_74_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08194_ net37 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07145_ _02301_ _02307_ _02585_ _02775_ _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_14_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07076_ _02658_ _02695_ _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06027_ _01682_ _01684_ _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_76_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07978_ ci_neuron.uut_simple_neuron.titan_id_2\[24\] ci_neuron.uut_simple_neuron.titan_id_5\[24\]
+ _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06929_ _02560_ _02563_ _02564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09717_ _00296_ net149 internal_ih.received_byte_count\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08503__A2 _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09648_ ci_neuron.stream_o\[25\] ci_neuron.output_memory\[25\] _04821_ _04823_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_84_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09579_ _04768_ _04782_ _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10285_ _00578_ net139 ci_neuron.stream_o\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04851__I1 internal_ih.byte3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08886__I _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout231_I net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05260_ _00908_ _00919_ _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05191_ _00865_ _00866_ _00868_ _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_3_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08950_ _04321_ _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07901_ _03481_ _03482_ _03483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09230__I0 _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08881_ _04282_ _00349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08733__A2 _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07832_ ci_neuron.uut_simple_neuron.titan_id_2\[1\] ci_neuron.uut_simple_neuron.titan_id_5\[1\]
+ _03424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_71_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07763_ _03364_ _03366_ _03367_ _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_79_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09502_ _03852_ ci_neuron.input_memory\[1\]\[19\] _01264_ _02552_ _04716_ _04717_
+ _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_04975_ _00681_ _00036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06714_ _02259_ _02298_ _02352_ _02353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07694_ ci_neuron.uut_simple_neuron.titan_id_4\[8\] ci_neuron.uut_simple_neuron.titan_id_3\[8\]
+ _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08497__A1 _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06645_ _02226_ _02231_ _02284_ _02285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09433_ _04652_ _04658_ _04659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09364_ _00727_ _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06576_ _01954_ _02192_ _02216_ _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09297__I0 _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08315_ ci_neuron.uut_simple_neuron.x0\[16\] _03823_ _03816_ _03818_ _03814_ _03830_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_05527_ _01172_ _01195_ _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09295_ ci_neuron.input_memory\[1\]\[8\] _04556_ _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05458_ _01084_ _01085_ _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08246_ _03769_ _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08177_ _03711_ _00085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07128_ _02716_ _02718_ _02759_ _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_05389_ _01035_ _01057_ _01060_ _01008_ _01061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_70_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07059_ _02184_ _02691_ _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06983__A1 _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05395__I _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10070_ _00197_ net200 ci_neuron.uut_simple_neuron.titan_id_0\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09221__I0 _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08488__A1 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10268_ _00561_ net152 ci_neuron.stream_o\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10199_ _00125_ net269 ci_neuron.uut_simple_neuron.titan_id_5\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06430_ _02038_ _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06361_ _01844_ _01902_ _02007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06292_ _01920_ _01924_ _01939_ _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_83_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05312_ _00968_ _00974_ _00985_ _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08100_ _03643_ _03645_ _03647_ _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09080_ _04389_ _04423_ _04424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05243_ _00909_ _00918_ _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08031_ _03589_ _00089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05174_ _00741_ _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09982_ _00497_ net109 ci_neuron.input_memory\[1\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout94_I net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ _04311_ _04312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_110_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08864_ internal_ih.byte1\[4\] internal_ih.byte0\[4\] _04270_ _04273_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07815_ _03411_ _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08795_ _04040_ _01098_ _04231_ _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07746_ _03352_ _03353_ _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04958_ internal_ih.byte0\[5\] _00670_ _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_84_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07677_ _03288_ _03293_ _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09416_ _04604_ _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_04889_ _00630_ _00012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06628_ _02266_ _02267_ _02268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_109_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06559_ _00163_ _02121_ _02153_ _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_63_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09347_ _04122_ ci_neuron.input_memory\[1\]\[31\] _04583_ _04587_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_51_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09278_ ci_neuron.input_memory\[1\]\[1\] _04546_ _04548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08229_ ci_neuron.uut_simple_neuron.x0\[7\] _03755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10122_ _00246_ net238 ci_neuron.uut_simple_neuron.titan_id_4\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10053_ _00538_ net165 ci_neuron.output_val_internal\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05930_ _01563_ _01589_ _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05861_ _00780_ _01469_ _01482_ _01522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_28_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07600_ _03216_ _03223_ _03224_ _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08580_ _03839_ _04049_ _04026_ _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07531_ _03106_ _03116_ _03156_ _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05792_ _01421_ _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07462_ _02937_ _03088_ _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06413_ _02057_ _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07393_ _03016_ _03020_ _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09201_ _03754_ _04500_ _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06344_ _01958_ _01968_ _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09132_ _04462_ _00420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08624__A1 _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06275_ _01899_ _01908_ _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09063_ _04383_ ci_neuron.stream_o\[3\] ci_neuron.stream_o\[19\] _04384_ _04407_
+ _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_05226_ _00878_ _00882_ _00902_ _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_4_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08014_ _03573_ _03574_ _03576_ _03577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05157_ ci_neuron.uut_simple_neuron.x2\[2\] ci_neuron.uut_simple_neuron.x2\[3\] ci_neuron.uut_simple_neuron.x2\[4\]
+ _00793_ _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_4_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05610__A1 _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05088_ _00760_ _00767_ _00769_ _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09965_ _00480_ net204 ci_neuron.input_memory\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08916_ _04302_ _00364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09896_ _00001_ net15 ci_neuron.address_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08847_ internal_ih.byte0\[5\] internal_ih.spi_rx_byte_i\[5\] _04258_ _04263_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08778_ _00867_ _04221_ _04223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07729_ _03339_ _00101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09256__S _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10105_ _00229_ net280 ci_neuron.uut_simple_neuron.titan_id_4\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10036_ _00521_ net169 ci_neuron.output_val_internal\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06060_ _01709_ _01716_ _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_53_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05011_ internal_ih.byte3\[4\] _00701_ _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_117_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06962_ _02538_ _02594_ _02595_ _02596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09750_ _00329_ net94 ci_neuron.uut_simple_neuron.x2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09681_ _00268_ net250 ci_neuron.uut_simple_neuron.x3\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05913_ _01532_ _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08701_ _04133_ _04162_ _04163_ _00288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06893_ _02484_ _02512_ _02527_ _02528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08632_ _03229_ _03941_ _04105_ _00277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05844_ _01403_ _01505_ _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08563_ _04047_ _00266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05775_ _00886_ _01178_ _01421_ _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_68_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07514_ _03068_ _03140_ _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08494_ _03753_ _03976_ _03755_ _03988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07445_ _02998_ _03039_ _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_81_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout15 net16 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout26 net27 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout37 ci_neuron.uut_simple_neuron.x0\[0\] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout59 net61 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout48 net49 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07376_ _03002_ _03003_ _03004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06327_ _01924_ _01939_ _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09115_ ci_neuron.uut_simple_neuron.titan_id_6\[1\] _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06258_ _01853_ _01906_ _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_60_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09046_ _04389_ _04392_ _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05209_ _00859_ _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06189_ _01821_ _01837_ _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09948_ _00463_ net107 ci_neuron.uut_simple_neuron.x0\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09879_ _00039_ net24 ci_neuron.value_i\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10019_ ci_neuron.input_memory\[1\]\[19\] net109 ci_neuron.uut_simple_neuron.titan_id_1\[21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout261_I net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05560_ _00749_ _01227_ _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_47_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05491_ _01078_ _01159_ _01160_ _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07230_ _02858_ _02859_ _02860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_119_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07161_ _02790_ _02758_ _02791_ _02792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__04864__A2 _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06112_ _01762_ _01767_ _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07092_ _02721_ _02722_ _02723_ _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06043_ _01661_ _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout205 net206 net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09555__A2 _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout238 net240 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout227 net231 net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout216 net217 net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09802_ _00381_ net53 internal_ih.byte6\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout249 net250 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07994_ ci_neuron.uut_simple_neuron.titan_id_2\[25\] ci_neuron.uut_simple_neuron.titan_id_5\[25\]
+ _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06945_ _02464_ _02463_ _02518_ _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09733_ _00312_ net228 ci_neuron.uut_simple_neuron.x2\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06876_ _02487_ _02511_ _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09664_ _00251_ net275 ci_neuron.uut_simple_neuron.x3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05827_ _01456_ _01488_ _01489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09595_ ci_neuron.stream_o\[2\] ci_neuron.output_memory\[2\] _04790_ _04793_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09423__I _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08615_ ci_neuron.value_i\[25\] _04032_ _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05758_ _01377_ _01419_ _01420_ _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08546_ ci_neuron.value_i\[14\] _04032_ _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05689_ _01316_ _01317_ _01352_ _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_49_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08477_ _03971_ _03972_ _03973_ _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_07428_ _02920_ _02972_ _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07359_ _02781_ _02834_ _02987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09029_ _04374_ _04376_ _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07557__A1 _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07309__A1 ci_neuron.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09537__A2 _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04991_ _00690_ _00043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06730_ _02364_ _02367_ _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06661_ _02244_ _02255_ _02300_ _02301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__09243__I _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05612_ _01235_ _01239_ _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08400_ _03903_ _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06592_ _02230_ _02232_ _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_52_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09380_ _00706_ ci_neuron.input_memory\[1\]\[1\] _00745_ _01848_ _04605_ _04607_
+ _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_05543_ _01011_ _01140_ _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_74_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08331_ _03836_ ci_neuron.uut_simple_neuron.x0\[20\] _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_19_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05474_ _01137_ _01143_ _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_74_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08262_ _03783_ _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_52_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07213_ _02779_ _02839_ _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08193_ ci_neuron.uut_simple_neuron.x0\[2\] _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_125_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07144_ _02701_ _02772_ _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_113_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07075_ _01889_ _02655_ _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06026_ _01594_ _01633_ _01683_ _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_76_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04850__I _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07977_ _03544_ _03545_ _03546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06928_ _02562_ _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09716_ _00295_ net148 internal_ih.received_byte_count\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06859_ _02384_ _02448_ _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09647_ _04822_ _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09578_ ci_neuron.uut_simple_neuron.x0\[31\] ci_neuron.input_memory\[1\]\[31\] ci_neuron.uut_simple_neuron.x2\[31\]
+ ci_neuron.uut_simple_neuron.x3\[31\] _04604_ _04606_ _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_38_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08529_ _04018_ _00261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_41_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10284_ _00577_ net141 ci_neuron.stream_o\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_49_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09542__I2 _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06269__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09207__A1 _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05190_ _00812_ _00846_ _00867_ _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_3_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07900_ ci_neuron.uut_simple_neuron.titan_id_2\[12\] ci_neuron.uut_simple_neuron.titan_id_5\[12\]
+ _03482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08880_ internal_ih.byte2\[3\] internal_ih.byte1\[3\] _04280_ _04282_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07831_ _03423_ _00138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_71_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_127_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07762_ ci_neuron.uut_simple_neuron.titan_id_4\[20\] ci_neuron.uut_simple_neuron.titan_id_3\[20\]
+ _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09501_ _04668_ _04717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04974_ internal_ih.byte1\[4\] _00680_ _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06713_ _02262_ _02297_ _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07693_ ci_neuron.uut_simple_neuron.titan_id_4\[8\] ci_neuron.uut_simple_neuron.titan_id_3\[8\]
+ ci_neuron.uut_simple_neuron.titan_id_4\[7\] ci_neuron.uut_simple_neuron.titan_id_3\[7\]
+ _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_94_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06644_ _02227_ _02283_ _02284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09432_ _03772_ ci_neuron.input_memory\[1\]\[9\] _00896_ _02089_ _04644_ _04645_
+ _04658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_06575_ _01955_ _02085_ _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_94_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05180__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09363_ _04597_ _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05526_ _01183_ _01194_ _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08314_ _03829_ _00177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09294_ _03990_ _04553_ _04557_ _00487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_25_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05457_ _01084_ _01085_ _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08245_ ci_neuron.uut_simple_neuron.x0\[8\] _03769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05388_ _01059_ _01060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08176_ _03709_ _03710_ _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_113_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07127_ _02720_ _02748_ _02758_ _02759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_104_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08421__A2 _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07058_ _02190_ _02690_ _02691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06009_ ci_neuron.uut_simple_neuron.x2\[28\] _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_89_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_43_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08799__I0 _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10144__D _00209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10267_ _00560_ net152 ci_neuron.stream_o\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10198_ _00124_ net269 ci_neuron.uut_simple_neuron.titan_id_5\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08479__A2 _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_109_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_61_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06360_ _01997_ _02005_ _02006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_84_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06291_ _01929_ _01935_ _01938_ _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_05311_ _00942_ _00984_ _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_126_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05242_ _00852_ _00912_ _00917_ _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_72_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08030_ ci_neuron.uut_simple_neuron.titan_id_1\[5\] ci_neuron.uut_simple_neuron.titan_id_0\[5\]
+ _03588_ _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_114_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05173_ _00806_ _00848_ _00849_ _00829_ _00850_ _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_12_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09981_ _00496_ net228 ci_neuron.input_memory\[1\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08932_ _04256_ _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__04976__A1 internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08863_ _04272_ _00341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07814_ ci_neuron.uut_simple_neuron.titan_id_4\[29\] ci_neuron.uut_simple_neuron.titan_id_3\[29\]
+ _03410_ _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08794_ _04232_ _00312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07745_ ci_neuron.uut_simple_neuron.titan_id_4\[18\] ci_neuron.uut_simple_neuron.titan_id_3\[18\]
+ _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04957_ _00671_ _00059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07676_ ci_neuron.uut_simple_neuron.titan_id_4\[6\] ci_neuron.uut_simple_neuron.titan_id_3\[6\]
+ _03295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04888_ internal_ih.byte4\[1\] _00625_ _00628_ internal_ih.byte0\[1\] _00630_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09415_ ci_neuron.output_memory\[7\] _04628_ _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06627_ _01921_ _02263_ _02264_ _02267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_75_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06558_ _02124_ _02152_ _02200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09346_ _04586_ _00510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_51_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04900__B2 internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04900__A1 internal_ih.byte4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06489_ _02098_ _02132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05509_ _01177_ _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_62_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09277_ _03947_ _04544_ _04547_ _00480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08228_ _03753_ _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08159_ ci_neuron.uut_simple_neuron.titan_id_1\[26\] ci_neuron.uut_simple_neuron.titan_id_0\[26\]
+ _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10121_ _00245_ net238 ci_neuron.uut_simple_neuron.titan_id_4\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04967__A1 internal_ih.byte1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10052_ _00537_ net165 ci_neuron.output_val_internal\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06708__A2 _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10139__D _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04958__A1 internal_ih.byte0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05860_ _00780_ _01469_ _01482_ _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09361__A3 _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05791_ _01415_ _01441_ _01452_ _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07530_ _03078_ _03104_ _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07461_ ci_neuron.uut_simple_neuron.x3\[27\] ci_neuron.uut_simple_neuron.x3\[28\]
+ _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07392_ _02812_ _03019_ _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06412_ _02055_ _02056_ _02057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09200_ _03979_ _04494_ _04501_ _00449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_17_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06343_ _01988_ _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09131_ ci_neuron.uut_simple_neuron.titan_id_6\[9\] _04462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09062_ _04405_ _04406_ _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06274_ _01898_ _01907_ _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05225_ _00879_ _00901_ _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08013_ ci_neuron.uut_simple_neuron.titan_id_2\[30\] ci_neuron.uut_simple_neuron.titan_id_5\[30\]
+ _03576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05156_ _00811_ ci_neuron.uut_simple_neuron.x2\[7\] _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05087_ _00760_ _00768_ _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09964_ _00479_ net122 spi_interface_cvonk.state\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08915_ internal_ih.byte4\[2\] internal_ih.byte3\[2\] _04301_ _04302_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09895_ _00057_ net19 ci_neuron.value_i\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05175__B _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08846_ _04262_ _00334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05989_ _01551_ _01642_ _01643_ _01646_ _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08777_ _03990_ _04218_ _04222_ _00305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07728_ ci_neuron.uut_simple_neuron.titan_id_4\[15\] ci_neuron.uut_simple_neuron.titan_id_3\[15\]
+ _03338_ _03339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_67_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07659_ ci_neuron.uut_simple_neuron.titan_id_4\[3\] ci_neuron.uut_simple_neuron.titan_id_3\[3\]
+ _03281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_48_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09329_ _04085_ ci_neuron.input_memory\[1\]\[23\] _04572_ _04577_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_106_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10104_ _00228_ net279 ci_neuron.uut_simple_neuron.titan_id_4\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08926__I0 internal_ih.byte4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10035_ _00520_ net169 ci_neuron.output_val_internal\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_106_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08606__A2 _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05010_ _00685_ _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_117_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06961_ _02540_ _02566_ _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09680_ _00267_ net232 ci_neuron.uut_simple_neuron.x3\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05912_ _01528_ _01569_ _01570_ _01571_ _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_08700_ internal_ih.spi_rx_byte_i\[6\] _04148_ _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06892_ _02487_ _02511_ _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08631_ _04011_ _04104_ _04105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05843_ _01497_ _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_89_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05774_ _01426_ _01432_ _01436_ _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_77_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08562_ _04046_ _02384_ _04028_ _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07513_ _03135_ _03139_ _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08493_ _03753_ _03755_ _03976_ _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_07444_ _03069_ _03070_ _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_81_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout38 ci_neuron.uut_simple_neuron.x2\[0\] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout27 net36 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout16 net17 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout49 net50 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07375_ _02942_ _02943_ _03003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06326_ _01924_ _01939_ _01973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09114_ _04453_ _00411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06257_ _01902_ _01905_ _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_60_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09045_ ci_neuron.output_val_internal\[25\] ci_neuron.output_val_internal\[17\] ci_neuron.output_val_internal\[9\]
+ ci_neuron.output_val_internal\[1\] _04390_ _04391_ _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_44_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05208_ _00841_ _00883_ _00884_ _00744_ _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06188_ _01821_ _01837_ _01840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_92_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05139_ _00744_ _00784_ _00798_ _00819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_8_Left_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09947_ _00462_ net100 ci_neuron.uut_simple_neuron.x0\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09878_ _00038_ net23 ci_neuron.value_i\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08829_ _04119_ _01793_ _04246_ _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05586__A1 _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08772__A1 _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10018_ ci_neuron.input_memory\[1\]\[18\] net110 ci_neuron.uut_simple_neuron.titan_id_1\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05490_ _01081_ _01113_ _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05510__A1 _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07160_ _02720_ _02748_ _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07263__A1 _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07091_ _02678_ _02684_ _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06111_ _01615_ _01766_ _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_124_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06042_ _01698_ _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout228 net230 net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout217 net291 net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout206 net207 net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09801_ _00380_ net54 internal_ih.byte6\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout239 net240 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09732_ _00311_ net228 ci_neuron.uut_simple_neuron.x2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07993_ _03546_ _03558_ _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06944_ _02411_ _02356_ _02410_ _02406_ _02467_ _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_06875_ _02491_ _02510_ _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09663_ _00250_ net264 ci_neuron.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05826_ _01460_ _01487_ _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08614_ _04090_ _00274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09594_ _04792_ _00552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08545_ _04000_ _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05757_ _01104_ _01188_ _01370_ _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_05688_ _01316_ _01317_ _01352_ _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09491__A2 _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08476_ ci_neuron.value_i\[4\] _03951_ _03973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07427_ _02996_ _03054_ _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_17_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09618__I1 ci_neuron.output_memory\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07358_ _02784_ _02833_ _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_116_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06309_ _01954_ _01955_ _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07289_ _02899_ _02907_ _02917_ _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_115_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09028_ _04191_ _04375_ _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09306__I0 _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07493__A1 _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09609__I1 ci_neuron.output_memory\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_62_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06599__A3 _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_114_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09671__D _00258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04990_ internal_ih.byte2\[3\] _00686_ _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_36_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06660_ _02258_ _02299_ _02300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05611_ _01248_ _01277_ _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_65_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06591_ _02142_ _02231_ _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_59_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05542_ _01018_ _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08330_ _03843_ _00179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05473_ _00864_ _01142_ _01143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08261_ ci_neuron.uut_simple_neuron.x0\[11\] _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07212_ _02842_ _00243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08192_ _03723_ _00066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07143_ _02771_ _02768_ _02772_ _02704_ _02773_ _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XPHY_EDGE_ROW_89_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07074_ _02706_ _00241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06025_ _01601_ _01632_ _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07976_ ci_neuron.uut_simple_neuron.titan_id_2\[25\] ci_neuron.uut_simple_neuron.titan_id_5\[25\]
+ _03545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06927_ _02279_ _02561_ _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_98_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09715_ _00294_ net148 internal_ih.received_byte_count\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09646_ ci_neuron.stream_o\[24\] ci_neuron.output_memory\[24\] _04821_ _04822_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06858_ _02447_ _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06789_ _01991_ _02375_ _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05809_ _00852_ _01469_ _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09577_ ci_neuron.output_memory\[31\] _04766_ _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08528_ _04017_ _02139_ _03969_ _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07475__A1 _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08459_ net37 ci_neuron.uut_simple_neuron.x0\[1\] ci_neuron.uut_simple_neuron.x0\[2\]
+ _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_108_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05789__A1 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10283_ _00576_ net141 ci_neuron.stream_o\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07950__A2 ci_neuron.uut_simple_neuron.titan_id_5\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09542__I3 _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout217_I net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07830_ _03421_ _03422_ _03423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07761_ ci_neuron.uut_simple_neuron.titan_id_4\[20\] ci_neuron.uut_simple_neuron.titan_id_3\[20\]
+ _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_127_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06712_ _02350_ _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09500_ _04666_ _04716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_04973_ _00664_ _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07692_ _03300_ _03305_ _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06643_ ci_neuron.uut_simple_neuron.x3\[14\] _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09431_ ci_neuron.output_memory\[9\] _04650_ _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06574_ _02177_ _02196_ _02214_ _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_fanout32_I net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09362_ _04596_ _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05525_ _01171_ _01193_ _01194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08313_ _03822_ _03824_ _03828_ _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_19_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09293_ ci_neuron.input_memory\[1\]\[7\] _04556_ _04557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05456_ _01082_ _01112_ _01125_ _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08244_ _03768_ _00198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05387_ _01058_ _01056_ _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_31_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08175_ ci_neuron.uut_simple_neuron.titan_id_1\[29\] ci_neuron.uut_simple_neuron.titan_id_0\[29\]
+ _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07126_ _02751_ _02757_ _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_112_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07057_ _02329_ _02628_ _02689_ _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06008_ _01621_ _01622_ _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_7_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07932__A2 ci_neuron.uut_simple_neuron.titan_id_5\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07959_ ci_neuron.uut_simple_neuron.titan_id_2\[22\] ci_neuron.uut_simple_neuron.titan_id_5\[22\]
+ _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09629_ _04812_ _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_26_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06120__A1 _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10266_ _00559_ net151 ci_neuron.stream_o\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10197_ _00123_ net269 ci_neuron.uut_simple_neuron.titan_id_5\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07439__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06290_ _01937_ _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05310_ _00868_ _00983_ _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05241_ _00913_ _00916_ _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05172_ _00831_ _00844_ _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09980_ _00495_ net112 ci_neuron.input_memory\[1\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08931_ _04310_ _00371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08862_ internal_ih.byte1\[3\] internal_ih.byte0\[3\] _04270_ _04272_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07813_ _03387_ _03388_ _03404_ _03409_ _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_4_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08793_ _04034_ _01052_ _04231_ _04232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07744_ _03350_ _03351_ _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04956_ internal_ih.byte0\[4\] _00670_ _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07675_ _03294_ _00122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06626_ _02265_ _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04887_ _00629_ _00001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09414_ _04627_ _04639_ _04641_ _04642_ _00522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_109_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09419__A2 _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06557_ _02170_ _02198_ _02199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_90_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09345_ _04119_ ci_neuron.input_memory\[1\]\[30\] _04583_ _04586_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_51_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06488_ _02088_ _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05508_ _01173_ _01176_ _01042_ _01177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06102__A1 _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09276_ ci_neuron.input_memory\[1\]\[0\] _04546_ _04547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05439_ _01049_ _01050_ _01048_ _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_63_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08227_ _03752_ _03753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_31_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08158_ ci_neuron.uut_simple_neuron.titan_id_1\[26\] ci_neuron.uut_simple_neuron.titan_id_0\[26\]
+ _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07109_ _02441_ _02740_ _02741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08089_ _03634_ _03636_ _03638_ _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10120_ _00244_ net239 ci_neuron.uut_simple_neuron.titan_id_4\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10051_ _00536_ net166 ci_neuron.output_val_internal\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05916__A1 _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_59_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05080__A1 _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10249_ _00146_ net101 ci_neuron.uut_simple_neuron.titan_id_6\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout284_I net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05907__A1 _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05790_ _01418_ _01440_ _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06580__A1 _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07460_ _03085_ _03086_ _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07391_ _03017_ _03018_ _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06411_ _01860_ _01931_ _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06342_ _01953_ _01988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09130_ _04461_ _00419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09061_ _04358_ ci_neuron.stream_o\[11\] _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06273_ _01894_ _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08012_ _03575_ _00150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05224_ _00885_ _00900_ _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05155_ _00832_ _00833_ _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05086_ _00766_ _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09963_ _00478_ net128 spi_interface_cvonk.state\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08914_ _04290_ _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09894_ _00056_ net19 ci_neuron.value_i\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08845_ internal_ih.byte0\[4\] internal_ih.spi_rx_byte_i\[4\] _04258_ _04262_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08776_ _00847_ _04221_ _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08560__A2 _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05988_ _01644_ _01645_ _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07727_ _03334_ _03335_ _03337_ _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09442__I _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04939_ internal_ih.byte6\[5\] _00658_ _00659_ internal_ih.byte2\[5\] _00661_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07658_ _03280_ _00118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07589_ _03145_ _03214_ _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06609_ _02209_ _02249_ _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09328_ _04079_ _04546_ _04576_ _00502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09259_ _04383_ _04373_ _04374_ _04533_ _00476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08871__I0 internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05210__I _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10103_ _00169_ net279 ci_neuron.uut_simple_neuron.titan_id_4\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09328__A1 _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10034_ _00519_ net144 ci_neuron.output_val_internal\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06865__A2 ci_neuron.uut_simple_neuron.x3\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08862__I0 internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09406__I2 _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09567__A1 ci_neuron.output_memory\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09674__D _00261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09527__I _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06960_ _02540_ _02566_ _02594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input4_I sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06891_ _02476_ _02483_ _02525_ _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05911_ _01527_ _01536_ _01571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08917__I1 internal_ih.byte3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05842_ _01408_ _01503_ _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08630_ _04101_ _04103_ _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06553__A1 _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05773_ _01425_ _01435_ _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08561_ _03996_ _04042_ _04044_ _04045_ _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_07512_ _03137_ _03138_ _03139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08492_ _03940_ _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07443_ _03041_ _03052_ _03070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06856__A2 _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout17 net18 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout28 net29 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout39 net40 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07374_ _02932_ _02941_ _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout9_I net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09113_ ci_neuron.uut_simple_neuron.titan_id_6\[0\] _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06325_ _01947_ _01971_ _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06256_ _01873_ _01904_ _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09044_ internal_ih.data_pointer\[1\] _04391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05207_ _00842_ _00871_ _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_41_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06187_ _01837_ _01838_ _01839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_13_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05138_ _00814_ _00817_ _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06792__A1 _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05069_ ci_neuron.uut_simple_neuron.x2\[2\] _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09946_ _00461_ net100 ci_neuron.uut_simple_neuron.x0\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09877_ _00037_ net32 ci_neuron.value_i\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06544__A1 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08828_ _04251_ _00327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08759_ _00737_ _04211_ _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_109_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09549__A1 ci_neuron.output_val_internal\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_118_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10017_ ci_neuron.input_memory\[1\]\[17\] net112 ci_neuron.uut_simple_neuron.titan_id_1\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_127_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout247_I net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_119_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07090_ _02686_ _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_82_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06110_ _01613_ _01765_ _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_124_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06041_ _01255_ _01697_ _01698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_124_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05785__I _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout218 net220 net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout229 net230 net229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout207 net213 net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09800_ _00379_ net48 internal_ih.byte6\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07992_ _03552_ _03554_ _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06943_ _02577_ _02521_ _02578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09731_ _00310_ net253 ci_neuron.uut_simple_neuron.x2\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07971__B1 _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06874_ _02493_ _02509_ _02510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09662_ _04830_ _00582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05825_ _01467_ _01486_ _01487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08613_ _04089_ _02865_ _04086_ _04090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09593_ ci_neuron.stream_o\[1\] ci_neuron.output_memory\[1\] _04790_ _04792_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05756_ _01333_ _01372_ _01145_ _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_08544_ _03808_ _04030_ _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05687_ _01236_ _01351_ _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08475_ _03739_ _03963_ _03972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07426_ _03040_ _03053_ _03054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_119_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09079__I0 ci_neuron.output_val_internal\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07357_ _02985_ _00245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06308_ _01933_ _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07288_ _02902_ _02906_ _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09027_ _04152_ _04172_ _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06239_ _01888_ _00166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__04863__I1 internal_ih.byte3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09929_ _00444_ net189 ci_neuron.uut_simple_neuron.x0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_103_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08690__A1 _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09490__I0 _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_114_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05008__A1 internal_ih.byte3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05610_ _01124_ _01276_ _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_129_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06590_ _02227_ ci_neuron.uut_simple_neuron.x3\[14\] _02231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05541_ _01180_ _01208_ _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05472_ _01139_ _01141_ _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08260_ _03776_ _03782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07211_ _02778_ _02841_ _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08808__I0 _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08191_ ci_neuron.uut_simple_neuron.titan_id_1\[2\] ci_neuron.uut_simple_neuron.titan_id_0\[2\]
+ _03723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07142_ _02647_ _02765_ _02764_ _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_54_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07236__A2 _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07073_ _02700_ _02705_ _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06024_ _01648_ _01681_ _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09233__I0 _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07975_ ci_neuron.uut_simple_neuron.titan_id_2\[25\] ci_neuron.uut_simple_neuron.titan_id_5\[25\]
+ _03544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06926_ _02232_ _02386_ _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09714_ _00293_ net148 internal_ih.received_byte_count\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06857_ _02452_ _02455_ _02492_ _02493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07235__I ci_neuron.uut_simple_neuron.x3\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09645_ _04810_ _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05808_ _01432_ _01436_ _01468_ _01469_ _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_69_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06788_ _01969_ _02374_ _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09576_ _04765_ _04777_ _04779_ _04780_ _00546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05739_ _01356_ _01402_ _01354_ _01403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08527_ _04013_ _04014_ _04015_ _04016_ _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_92_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08458_ _03940_ _03957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07409_ _03034_ _03036_ _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08389_ _03886_ _03887_ _03895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09224__I0 _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10282_ _00575_ net141 ci_neuron.stream_o\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06910__A1 _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09679__CLK net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08415__A1 _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06977__A1 _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09215__I0 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07760_ _03365_ _00106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04972_ _00679_ _00035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_127_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06711_ _02266_ _02311_ _02349_ _02350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07691_ _03287_ _03296_ _03307_ _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09430_ _04649_ _04651_ _04654_ _04656_ _00524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06642_ _02136_ _02233_ _02281_ _02282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06573_ _02180_ _02195_ _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09361_ _04595_ _00724_ _03923_ _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_129_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05524_ _01147_ _01188_ _01189_ _01192_ _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_09292_ _04545_ _04556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08312_ _03826_ _03827_ _03828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08243_ _03766_ _03767_ _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_117_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05455_ _01108_ _01111_ _01125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05386_ _00741_ _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08174_ _03704_ _03705_ _03708_ _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07125_ _02754_ _02756_ _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07056_ _02330_ _02494_ _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_70_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06007_ _01662_ _01664_ _01665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09445__I _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07958_ _03520_ _03525_ _03526_ _03528_ _03529_ _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_06909_ _02131_ _02543_ _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_69_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07889_ _03467_ _03468_ _03469_ _03471_ _03472_ _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_97_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09628_ ci_neuron.stream_o\[16\] ci_neuron.output_memory\[16\] _04811_ _04812_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_26_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09559_ _00727_ _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_54_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05459__A1 _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06959__A1 _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10265_ _00558_ net153 ci_neuron.stream_o\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10196_ _00122_ net269 ci_neuron.uut_simple_neuron.titan_id_5\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_70_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_122_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05240_ _00914_ _00915_ _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05171_ _00831_ _00844_ _00849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_25_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06889__I _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05622__A1 _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08930_ internal_ih.byte5\[1\] internal_ih.byte4\[1\] _04306_ _04310_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08861_ _04271_ _00340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07812_ ci_neuron.uut_simple_neuron.titan_id_4\[28\] ci_neuron.uut_simple_neuron.titan_id_3\[28\]
+ _03403_ _03406_ _03408_ _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_4_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08792_ _04224_ _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07743_ _03347_ _03348_ _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04955_ _00664_ _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07674_ _03292_ _03293_ _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04886_ internal_ih.byte4\[0\] _00625_ _00628_ internal_ih.byte0\[0\] _00629_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06625_ _02263_ _02264_ _01921_ _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09413_ ci_neuron.output_val_internal\[6\] _04633_ _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06556_ _02172_ _02197_ _02198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09344_ _04585_ _00509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_51_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06487_ _01850_ _02129_ _02130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05507_ _00981_ _01140_ _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_62_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09275_ _04545_ _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05438_ _01049_ _01048_ _01050_ _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08226_ ci_neuron.uut_simple_neuron.x0\[6\] _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05861__A1 _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08157_ _03694_ _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07108_ _02390_ _02615_ _02740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05369_ _01013_ _01014_ _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08088_ ci_neuron.uut_simple_neuron.titan_id_1\[13\] ci_neuron.uut_simple_neuron.titan_id_0\[13\]
+ _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07039_ _02619_ _02627_ _02672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10050_ _00535_ net136 ci_neuron.output_val_internal\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08618__A1 _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09291__A1 _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10248_ _00145_ net81 ci_neuron.uut_simple_neuron.titan_id_6\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10179_ _00076_ net108 ci_neuron.uut_simple_neuron.titan_id_2\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06410_ _01858_ _02055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07390_ _02676_ _02858_ _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_17_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06341_ _01985_ _01986_ _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09282__A1 _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06272_ _01891_ _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06096__A1 _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09060_ _04360_ _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05223_ _00889_ _00899_ _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08880__I1 internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08011_ _03573_ _03574_ _03575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05154_ ci_neuron.uut_simple_neuron.x2\[2\] ci_neuron.uut_simple_neuron.x2\[3\] ci_neuron.uut_simple_neuron.x2\[4\]
+ ci_neuron.uut_simple_neuron.x2\[5\] _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_12_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05085_ _00756_ _00766_ _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09962_ _00477_ net122 spi_interface_cvonk.state\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08913_ _04300_ _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09893_ _00054_ net19 ci_neuron.value_i\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08844_ _04261_ _00333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05987_ _01634_ _01636_ _01638_ _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08775_ _04210_ _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07726_ ci_neuron.uut_simple_neuron.titan_id_4\[14\] ci_neuron.uut_simple_neuron.titan_id_3\[14\]
+ _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_04938_ _00660_ _00013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07657_ ci_neuron.uut_simple_neuron.titan_id_4\[3\] ci_neuron.uut_simple_neuron.titan_id_3\[3\]
+ _03279_ _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_04869_ _00605_ _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_36_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07588_ _03146_ _03213_ _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06608_ _02244_ _02248_ _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06539_ _02141_ _02181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09327_ ci_neuron.input_memory\[1\]\[22\] _04556_ _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08871__I1 internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09258_ _04381_ _04384_ _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09189_ _04488_ _04494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08209_ _03733_ _03737_ _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08802__I _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10102_ _00168_ net276 ci_neuron.uut_simple_neuron.titan_id_4\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09328__A2 _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06322__I _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10033_ _00518_ net144 ci_neuron.output_val_internal\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08000__A2 ci_neuron.uut_simple_neuron.titan_id_5\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09406__I3 _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06890_ _02479_ _02482_ _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05910_ _01530_ _01534_ _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05841_ _01450_ _01443_ _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05772_ _01430_ _01434_ _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08560_ ci_neuron.value_i\[16\] _04001_ _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07511_ _02993_ _03055_ _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08491_ _03957_ _03984_ _03985_ _00256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07442_ _03042_ _03043_ _03051_ _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout18 net27 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout29 net30 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_33_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07373_ _02945_ _02948_ _03000_ _03001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04867__A2 _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06324_ _01951_ _01970_ _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09112_ _04415_ _04451_ _04452_ _00410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06255_ ci_neuron.uut_simple_neuron.x3\[5\] _01903_ _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09043_ internal_ih.data_pointer\[0\] _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06186_ ci_neuron.uut_simple_neuron.x3\[3\] _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05206_ _00853_ _00871_ _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05137_ _00781_ _00816_ _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07238__I ci_neuron.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06241__A1 _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05068_ _00737_ _00751_ _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09945_ _00460_ net104 ci_neuron.uut_simple_neuron.x0\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09876_ _00036_ net32 ci_neuron.value_i\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08827_ _04116_ _01751_ _04246_ _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08758_ _04210_ _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07709_ _03323_ _00097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08689_ internal_ih.spi_rx_byte_i\[3\] _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09494__A1 ci_neuron.output_memory\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08541__I0 _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10016_ ci_neuron.input_memory\[1\]\[16\] net112 ci_neuron.uut_simple_neuron.titan_id_1\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_19_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__04849__A2 _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09237__A1 _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_119_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06040_ _01179_ _01696_ _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_78_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout219 net220 net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout208 net209 net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07991_ _03557_ _00146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06942_ _02463_ _02465_ _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09730_ _00309_ net254 ci_neuron.uut_simple_neuron.x2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06873_ _02505_ _02508_ _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09661_ ci_neuron.stream_o\[31\] ci_neuron.output_memory\[31\] _04826_ _04830_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05824_ _01470_ _01485_ _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09592_ _04791_ _00551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08612_ ci_neuron.value_i\[24\] _04088_ _03953_ _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05755_ _01416_ _01387_ _01417_ _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08543_ _03794_ _03796_ _04015_ _04030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_49_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05686_ _01319_ _01350_ _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08474_ _03942_ _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_07425_ _03041_ _03052_ _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_64_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07356_ _02979_ _02984_ _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07287_ _02910_ _02912_ _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06307_ _01931_ _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06238_ _01885_ _01887_ _01888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09026_ _04145_ _04179_ _04373_ _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06169_ _01820_ _01822_ _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06214__A1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09928_ _00443_ net130 internal_ih.received_byte_count\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09183__I _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09554__I2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09859_ _00438_ net68 ci_neuron.output_memory\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08262__I _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05540_ _00961_ _01207_ _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_129_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05471_ _00982_ _01017_ _01140_ _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07210_ _02840_ _02841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08190_ _03722_ _00087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07141_ _02700_ _02764_ _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_82_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07072_ _02587_ _02701_ _02704_ _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_124_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06023_ _01652_ _01680_ _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06747__A2 _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07516__I _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07974_ _03543_ _00143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06925_ _02550_ _02559_ _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09536__I2 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09713_ _00292_ net129 internal_ih.received_byte_count\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06856_ _02444_ _02451_ _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09644_ _04820_ _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05807_ _01435_ _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06787_ _02369_ _02399_ _02423_ _02424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09575_ ci_neuron.output_val_internal\[30\] _04771_ _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05738_ _01353_ _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08526_ ci_neuron.value_i\[11\] _03965_ _04016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05669_ ci_neuron.uut_simple_neuron.x2\[19\] ci_neuron.uut_simple_neuron.x2\[20\]
+ _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08457_ _03941_ _03955_ _03956_ _00251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_41_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07408_ _02041_ _03035_ _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08388_ _03893_ _03889_ _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07339_ _01929_ _02420_ _02317_ _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_61_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08082__I _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09009_ internal_ih.data_pointer\[1\] _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10281_ _00574_ net155 ci_neuron.stream_o\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06330__I _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06910__A2 _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04921__B2 internal_ih.byte1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout105_I net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06240__I _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04971_ internal_ih.byte1\[3\] _00675_ _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_127_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06710_ _02319_ _02348_ _02349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_79_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07690_ _03295_ _03298_ _03307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06641_ _02279_ _02280_ _02281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_78_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06572_ _01827_ _02212_ _02213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09360_ _00708_ _00729_ _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05523_ _01190_ _01191_ _01186_ _01192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_75_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09291_ _03984_ _04553_ _04555_ _00486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08311_ _03814_ _03819_ _03827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05454_ _00934_ _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_86_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08242_ _03765_ _03761_ _03764_ _03767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_7_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout18_I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05385_ _01056_ _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08173_ _03707_ _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07124_ _01882_ _02755_ _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08831__S _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07055_ _02675_ _02687_ _02688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_70_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06006_ _01663_ _01624_ _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07957_ ci_neuron.uut_simple_neuron.titan_id_2\[21\] ci_neuron.uut_simple_neuron.titan_id_5\[21\]
+ _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06908_ _02098_ _02542_ _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07888_ ci_neuron.uut_simple_neuron.titan_id_2\[9\] ci_neuron.uut_simple_neuron.titan_id_5\[9\]
+ _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06839_ _01984_ _02009_ _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09627_ _04810_ _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_26_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09558_ _04696_ _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08509_ _04000_ _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_108_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09489_ ci_neuron.output_memory\[17\] _04698_ _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_92_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08805__I _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Left_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08540__I _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10264_ _00557_ net184 ci_neuron.stream_o\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10195_ _00121_ net267 ci_neuron.uut_simple_neuron.titan_id_5\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09371__I _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_109_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05404__I _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08636__A2 _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_126_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05170_ _00814_ _00847_ _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_4_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07072__A1 _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08860_ internal_ih.byte1\[2\] internal_ih.byte0\[2\] _04270_ _04271_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07811_ _03407_ _03408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08791_ _04230_ _00311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07742_ ci_neuron.uut_simple_neuron.titan_id_4\[17\] ci_neuron.uut_simple_neuron.titan_id_3\[17\]
+ _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_79_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04954_ _00669_ _00058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05138__A1 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07673_ ci_neuron.uut_simple_neuron.titan_id_4\[6\] ci_neuron.uut_simple_neuron.titan_id_3\[6\]
+ _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04885_ _00627_ _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06624_ _01871_ _02218_ _02264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09412_ _04630_ _04640_ _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09343_ _04116_ ci_neuron.input_memory\[1\]\[29\] _04583_ _04585_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06555_ _02177_ _02196_ _02197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_90_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_51_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08627__A2 _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06486_ _02125_ _02128_ _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05506_ _00887_ _01142_ _01174_ _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_75_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09274_ _04542_ _04545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05437_ _01088_ _01095_ _01107_ _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08225_ _03751_ _00196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_99_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05368_ _01013_ _01014_ _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_31_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08156_ _03692_ _03693_ _03694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07107_ _02729_ _02738_ _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05299_ _00971_ _00972_ _00965_ _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08087_ _03637_ _00068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07038_ _02612_ _02669_ _02670_ _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08989_ internal_ih.current_instruction\[2\] _04341_ _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_39_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10247_ _00144_ net98 ci_neuron.uut_simple_neuron.titan_id_6\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08554__A1 _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10178_ _00075_ net110 ci_neuron.uut_simple_neuron.titan_id_2\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05540__A1 _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09657__I1 ci_neuron.output_memory\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06340_ _01830_ _01877_ _01892_ _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06271_ _01890_ _01917_ _01918_ _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06096__A2 _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05222_ _00890_ _00898_ _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_71_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08010_ ci_neuron.uut_simple_neuron.titan_id_2\[30\] ci_neuron.uut_simple_neuron.titan_id_5\[30\]
+ _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05153_ _00787_ _00816_ _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05084_ ci_neuron.uut_simple_neuron.x2\[4\] _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09961_ _00476_ net141 internal_ih.data_pointer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08912_ internal_ih.byte4\[1\] internal_ih.byte3\[1\] _04296_ _04300_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_110_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09892_ _00053_ net21 ci_neuron.value_i\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08843_ internal_ih.byte0\[3\] _04155_ _04258_ _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05986_ _01634_ _01636_ _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08774_ _03984_ _04218_ _04220_ _00304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07725_ _03336_ _00100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09345__I0 _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04937_ internal_ih.byte6\[4\] _00658_ _00659_ internal_ih.byte2\[4\] _00660_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06859__A1 _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06323__A3 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ _03275_ _03277_ _03278_ _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_04868_ _00615_ _00028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_36_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07587_ _03150_ _03212_ _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06607_ _02246_ _02247_ _02248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09648__I1 ci_neuron.output_memory\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06538_ _02147_ _02149_ _02179_ _02180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09326_ _04575_ _00501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09257_ _04532_ _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06469_ _02030_ _02016_ _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08208_ _03734_ _03735_ _03736_ _03737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09025__A2 _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09188_ _03955_ _04489_ _04493_ _00445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08139_ _03676_ _03678_ _03679_ _03680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_120_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10101_ _00167_ net274 ci_neuron.uut_simple_neuron.titan_id_4\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10032_ _00517_ net155 ci_neuron.output_val_internal\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07434__I _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09336__I0 _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_106_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09639__I1 ci_neuron.output_memory\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05589__A1 _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08527__A1 _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05840_ _01307_ _01312_ _01501_ _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_55_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07510_ _03136_ _03054_ _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05771_ _01433_ _01380_ _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_89_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08490_ _01959_ _03980_ _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07441_ _03067_ _03058_ _03068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_119_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05513__A1 _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout19 net22 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_33_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07372_ _02999_ _02944_ _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06323_ _01953_ _01958_ _01969_ _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09111_ internal_ih.spi_tx_byte_o\[7\] _04427_ _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06254_ ci_neuron.uut_simple_neuron.x3\[6\] _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09042_ _04355_ _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06185_ ci_neuron.uut_simple_neuron.x3\[2\] _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05205_ _00879_ _00873_ _00881_ _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_4_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05136_ _00794_ _00796_ _00815_ _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_40_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05067_ _00750_ _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09944_ _00459_ net114 ci_neuron.uut_simple_neuron.x0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05044__A3 _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08518__A1 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09875_ _00035_ net32 ci_neuron.value_i\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08826_ _04250_ _00326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09191__A1 _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09318__I0 _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05969_ _01609_ _01627_ _01628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08757_ _04207_ _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07708_ ci_neuron.uut_simple_neuron.titan_id_4\[11\] ci_neuron.uut_simple_neuron.titan_id_3\[11\]
+ _03322_ _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08688_ internal_ih.spi_tx_byte_o\[2\] _04137_ _04142_ _04152_ _04154_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07639_ _03187_ _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08541__I1 _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07257__A1 _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09309_ _04565_ _00494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_101_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10015_ ci_neuron.input_memory\[1\]\[15\] net113 ci_neuron.uut_simple_neuron.titan_id_1\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09237__A2 _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_78_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout209 net212 net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07990_ _03554_ _03556_ _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06941_ _02573_ _02575_ _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07971__A2 ci_neuron.uut_simple_neuron.titan_id_5\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09660_ _04829_ _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07074__I _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06872_ _02507_ _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08611_ _03877_ _03869_ _04077_ _04088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05734__A1 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05823_ _01471_ _01482_ _01484_ _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09591_ ci_neuron.stream_o\[0\] ci_neuron.output_memory\[0\] _04790_ _04791_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08542_ _04029_ _00263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05754_ _01388_ _01392_ _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07487__A1 _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08473_ _03970_ _00253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_46_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07424_ _03044_ _03051_ _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_119_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05685_ _01284_ _01349_ _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_59_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08834__S _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07355_ _02778_ _02980_ _02983_ _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07239__A1 ci_neuron.uut_simple_neuron.x3\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07286_ _02915_ _00244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06306_ _01834_ _01952_ _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06237_ _01857_ _01864_ _01886_ _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09025_ _04178_ _00600_ _04186_ _04373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06168_ _01821_ _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05119_ _00786_ _00789_ _00799_ _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06099_ _01754_ _01667_ ci_neuron.uut_simple_neuron.x2\[30\] _01755_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_EDGE_ROW_68_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09927_ _00032_ net9 ci_neuron.instruction_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07962__A2 ci_neuron.uut_simple_neuron.titan_id_5\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09554__I3 _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09858_ _00437_ net63 ci_neuron.output_memory\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08809_ _04241_ _00318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09789_ _00368_ net43 internal_ih.byte4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09467__A2 _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07402__A1 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07953__A2 ci_neuron.uut_simple_neuron.titan_id_5\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05407__I _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05192__A2 _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout252_I net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05470_ _01091_ _01099_ _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07140_ _02647_ _02765_ _02764_ _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_125_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06682__B _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07071_ _02637_ _02702_ _02641_ _02703_ _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_30_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06022_ _01650_ _01679_ _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07944__A2 ci_neuron.uut_simple_neuron.titan_id_5\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09712_ _00291_ net129 internal_ih.received_byte_count\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07973_ _03541_ _03542_ _03543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06924_ _02442_ _02558_ _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__09536__I3 _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06855_ _02081_ _02490_ _02491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_93_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09643_ ci_neuron.stream_o\[23\] ci_neuron.output_memory\[23\] _04816_ _04820_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05806_ _01058_ _01384_ _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09574_ _04768_ _04778_ _04779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06786_ _02372_ _02398_ _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08525_ _03785_ _04006_ _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05737_ _01304_ _01355_ _01401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06132__A1 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05668_ _01185_ _01187_ _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08456_ _01848_ _03948_ _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05052__I _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07407_ _02436_ _02454_ _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08387_ _03875_ _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07338_ _01946_ _01989_ _01991_ _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_116_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05599_ ci_neuron.uut_simple_neuron.x2\[18\] _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_9_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07269_ _02898_ _01848_ _02713_ _02313_ _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XPHY_EDGE_ROW_76_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09008_ _04355_ _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10280_ _00573_ net155 ci_neuron.stream_o\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06199__B2 _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_85_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_29_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08538__I _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05897__I _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09369__I _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07926__A2 ci_neuron.uut_simple_neuron.titan_id_5\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_04970_ _00678_ _00034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10190__D ci_neuron.uut_simple_neuron.titan_id_3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06640_ _02232_ _02280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06571_ _02210_ _02211_ _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_86_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05522_ ci_neuron.uut_simple_neuron.x2\[15\] ci_neuron.uut_simple_neuron.x2\[16\]
+ ci_neuron.uut_simple_neuron.x2\[17\] _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_09290_ ci_neuron.input_memory\[1\]\[6\] _04549_ _04555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09300__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08310_ _03825_ _03821_ _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05453_ _01117_ _01120_ _01122_ _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08241_ _03761_ _03764_ _03765_ _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05384_ _00940_ _01055_ _01056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08172_ ci_neuron.uut_simple_neuron.titan_id_1\[28\] ci_neuron.uut_simple_neuron.titan_id_0\[28\]
+ _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07614__A1 ci_neuron.uut_simple_neuron.x3\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07123_ _02217_ _02237_ _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07054_ _02678_ _02684_ _02686_ _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_70_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06005_ _01616_ _01663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08590__A2 _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07956_ _03512_ _03513_ _03527_ _03528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06907_ _02222_ _02506_ _02541_ _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_98_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07887_ _03457_ _03458_ _03470_ _03471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06838_ _02431_ _02458_ _02473_ _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09626_ _03926_ _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06769_ _02351_ _02353_ _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_26_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09557_ _04743_ _04759_ _04763_ _04764_ _00543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_77_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09488_ _04697_ _04699_ _04703_ _04706_ _00532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08508_ _03950_ _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08439_ _03939_ _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08653__I0 _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10263_ _00556_ net183 ci_neuron.stream_o\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10194_ _00120_ net267 ci_neuron.uut_simple_neuron.titan_id_5\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout215_I net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05083__A1 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08947__I1 internal_ih.byte5\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07810_ ci_neuron.uut_simple_neuron.titan_id_4\[28\] ci_neuron.uut_simple_neuron.titan_id_3\[28\]
+ ci_neuron.uut_simple_neuron.titan_id_4\[27\] ci_neuron.uut_simple_neuron.titan_id_3\[27\]
+ _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08790_ _04027_ _01006_ _04225_ _04230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07741_ _03349_ _00103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04953_ internal_ih.byte0\[3\] _00665_ _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07672_ _03290_ _03291_ _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04884_ _00626_ _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06623_ _01883_ _02217_ _02263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09411_ _03754_ ci_neuron.input_memory\[1\]\[6\] _00814_ _01959_ _04622_ _04623_
+ _04640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_06554_ _02180_ _02195_ _02196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_87_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09342_ _04584_ _00508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout30_I net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05505_ _01042_ _01173_ _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_75_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06485_ _02127_ _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09273_ _04543_ _04544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09380__S0 _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05436_ _01059_ _01106_ _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08224_ _03747_ _03750_ _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_16_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05367_ _00976_ _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10095__D ci_neuron.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08155_ ci_neuron.uut_simple_neuron.titan_id_1\[26\] ci_neuron.uut_simple_neuron.titan_id_0\[26\]
+ _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07106_ _02617_ _02737_ _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05298_ _00971_ _00964_ _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08086_ _03634_ _03636_ _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07037_ _02614_ _02630_ _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09472__I _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08988_ _04343_ _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_3_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07939_ _03512_ _03513_ _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05129__A2 _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09609_ ci_neuron.stream_o\[8\] ci_neuron.output_memory\[8\] _04800_ _04801_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04888__A1 internal_ih.byte4\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06629__A2 _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09418__I2 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10246_ _00143_ net98 ci_neuron.uut_simple_neuron.titan_id_6\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10177_ _00074_ net112 ci_neuron.uut_simple_neuron.titan_id_2\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06270_ _01909_ _01911_ _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08490__A1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05221_ _00894_ _00897_ _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_72_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05152_ _00784_ _00821_ _00823_ _00810_ _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_69_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05083_ _00749_ _00754_ _00764_ _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_12_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09960_ _00475_ net82 ci_neuron.uut_simple_neuron.x0\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08911_ _04299_ _00362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09891_ _00052_ net20 ci_neuron.value_i\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08842_ _04170_ _04254_ _04260_ _00332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09593__I1 ci_neuron.output_memory\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05985_ _01492_ _01547_ _01548_ _01641_ _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08773_ _00814_ _04214_ _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07724_ _03334_ _03335_ _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04936_ _00626_ _00659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07655_ ci_neuron.uut_simple_neuron.titan_id_4\[2\] ci_neuron.uut_simple_neuron.titan_id_3\[2\]
+ _03278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06606_ _02204_ _02203_ _02247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_94_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04867_ internal_ih.byte7\[3\] _00606_ _00614_ _00610_ _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_36_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07586_ _03152_ _03211_ _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_87_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06537_ _02178_ _02146_ _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09325_ _04074_ ci_neuron.input_memory\[1\]\[21\] _04572_ _04575_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08856__I0 internal_ih.byte1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06468_ _02073_ _02108_ _02111_ _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_106_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09256_ _04122_ ci_neuron.uut_simple_neuron.x0\[31\] _04490_ _04532_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05419_ _01018_ _01046_ _01089_ _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08207_ ci_neuron.uut_simple_neuron.x0\[1\] ci_neuron.uut_simple_neuron.x0\[2\] _03736_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06399_ _02000_ _02044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09187_ _00706_ _04491_ _04493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08138_ ci_neuron.uut_simple_neuron.titan_id_1\[22\] ci_neuron.uut_simple_neuron.titan_id_0\[22\]
+ _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08069_ _03618_ _03619_ _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10100_ _00166_ net276 ci_neuron.uut_simple_neuron.titan_id_4\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10031_ _00516_ net143 ci_neuron.output_val_internal\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09336__I1 ci_neuron.input_memory\[1\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08847__I0 internal_ih.byte0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05286__B2 _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10229_ _00156_ net195 ci_neuron.uut_simple_neuron.titan_id_6\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout282_I net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05770_ ci_neuron.uut_simple_neuron.x2\[23\] _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07440_ _02993_ _03055_ _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07371_ _02926_ _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06322_ _01968_ _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09110_ ci_neuron.stream_o\[31\] _04416_ _04450_ _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08463__A1 _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09041_ _04383_ ci_neuron.stream_o\[1\] ci_neuron.stream_o\[17\] _04384_ _04387_
+ _04388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_06253_ _01872_ _01879_ _01901_ _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06184_ _01835_ _01836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_96_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05204_ _00818_ _00880_ _00872_ _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08215__A1 _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05135_ _00753_ _00793_ _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_41_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05066_ _00749_ _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09943_ _00458_ net114 ci_neuron.uut_simple_neuron.x0\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09874_ _00034_ net32 ci_neuron.value_i\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08825_ _04110_ _01792_ _04246_ _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05968_ _01526_ _01626_ _01627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05055__I _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08756_ _04208_ _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05899_ _01557_ _01541_ _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07707_ _03312_ _03318_ _03321_ _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_67_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08687_ _04134_ _04151_ _04153_ _00284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04919_ internal_ih.byte5\[5\] _00646_ _00647_ internal_ih.byte1\[5\] _00649_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07638_ _03261_ _03262_ _03263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07569_ _03126_ _03128_ _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08829__I0 _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09308_ _04034_ ci_neuron.input_memory\[1\]\[14\] _04561_ _04565_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08454__A1 ci_neuron.value_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09239_ _04085_ _03864_ _04519_ _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04866__I1 internal_ih.byte3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09254__I0 _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10014_ ci_neuron.input_memory\[1\]\[14\] net113 ci_neuron.uut_simple_neuron.titan_id_1\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_19_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_67_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08693__B2 _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_78_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06940_ _02519_ _02518_ _02574_ _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_91_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_105_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06871_ _02222_ _02506_ _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input2_I spi_cs_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05822_ _01428_ _01429_ _01483_ _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08610_ _04087_ _00273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09590_ _04789_ _04790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05753_ _01369_ _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08541_ _04027_ _02228_ _04028_ _04029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05684_ _01323_ _01348_ _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08472_ _03967_ _01872_ _03969_ _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07423_ _01892_ _03050_ _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08684__B2 _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_114_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07354_ _02981_ _02843_ _02982_ _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08914__I _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07285_ _02845_ _02914_ _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_127_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06305_ _01829_ _01876_ _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06236_ _01836_ _01839_ _01865_ _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09024_ ci_neuron.stream_o\[24\] _04354_ _04371_ _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06167_ ci_neuron.uut_simple_neuron.x3\[1\] _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05118_ _00790_ _00798_ _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06098_ ci_neuron.uut_simple_neuron.x2\[27\] _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_123_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05049_ _00733_ _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09926_ _00031_ net9 ci_neuron.instruction_i\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07175__A1 _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09857_ _00436_ net64 ci_neuron.output_memory\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08808_ _04069_ ci_neuron.uut_simple_neuron.x2\[20\] _04239_ _04241_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09788_ _00367_ net39 internal_ih.byte4\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08739_ _04193_ _04196_ _04197_ _00292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_103_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09490__I3 _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09390__I _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07070_ _02644_ _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_125_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07641__A2 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06021_ _01654_ _01678_ _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09711_ _00290_ net121 spi_interface_cvonk.buffer\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07972_ ci_neuron.uut_simple_neuron.titan_id_2\[24\] ci_neuron.uut_simple_neuron.titan_id_5\[24\]
+ _03542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06923_ _02554_ _02557_ _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06854_ _02053_ _02489_ _02490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09642_ _04819_ _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06785_ _02419_ _02421_ _02422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05805_ _01208_ _01389_ _01466_ _01467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09573_ _03916_ ci_neuron.input_memory\[1\]\[30\] _01793_ ci_neuron.uut_simple_neuron.x3\[30\]
+ _04760_ _04761_ _04778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_05736_ _01396_ _01399_ _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_77_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08524_ _04005_ _03998_ _03783_ _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05667_ _01186_ _01287_ _01223_ _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08455_ _00065_ _03952_ _03954_ _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07406_ _03032_ _03033_ _03034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05598_ _01227_ _01264_ _01265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08386_ _03891_ _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07337_ _02964_ _02965_ _02966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07268_ _01847_ _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_104_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07199_ _02827_ _02829_ _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06219_ _01858_ _01868_ _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_104_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09007_ _04177_ _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09909_ _00005_ net7 ci_neuron.address_i\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_29_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05634__A1 _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06570_ _01889_ _02176_ _02211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_86_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05521_ _01097_ _01149_ _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09300__A2 _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05452_ _01074_ _01077_ _01115_ _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_74_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08240_ ci_neuron.uut_simple_neuron.x0\[7\] ci_neuron.uut_simple_neuron.x0\[8\] _03765_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_117_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05873__A1 _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08171_ _03706_ _00084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07122_ _02752_ _02753_ _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05383_ _01053_ _01054_ _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07614__A2 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07053_ _02379_ _02685_ _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06004_ _01617_ _01623_ _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06050__A1 _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07955_ ci_neuron.uut_simple_neuron.titan_id_2\[19\] ci_neuron.uut_simple_neuron.titan_id_5\[19\]
+ _03527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06906_ _02223_ _02379_ _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07145__A4 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07886_ _03453_ _03460_ _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09625_ _04809_ _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06837_ _02434_ _02457_ _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06353__A2 _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06768_ _02405_ _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_26_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09556_ ci_neuron.output_val_internal\[27\] _04749_ _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06699_ ci_neuron.uut_simple_neuron.x3\[15\] ci_neuron.uut_simple_neuron.x3\[16\]
+ _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05719_ _01344_ _01328_ _01382_ _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_54_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08507_ _03770_ _03987_ _03772_ _03999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09487_ ci_neuron.output_val_internal\[16\] _04705_ _04706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08438_ _03938_ _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08369_ _03874_ _03877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10262_ _00555_ net155 ci_neuron.stream_o\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10193_ _00118_ net197 ci_neuron.uut_simple_neuron.titan_id_5\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06041__A1 _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06344__A2 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07541__A1 _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09294__A1 _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07740_ _03347_ _03348_ _03349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04952_ _00668_ _00055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_88_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07671_ _03287_ _03288_ _03291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04883_ _00603_ _00596_ _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06622_ _02213_ _02260_ _02261_ _02262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09410_ ci_neuron.output_memory\[6\] _04628_ _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06553_ _02191_ _02194_ _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09341_ _04110_ ci_neuron.input_memory\[1\]\[28\] _04583_ _04584_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05504_ _00981_ _01140_ _01173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06484_ _01896_ _01994_ _02126_ _02127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09272_ _04542_ _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09380__S1 _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05435_ _01098_ _01105_ _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08223_ _03748_ _03749_ _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_99_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05366_ _00972_ _01035_ _01037_ _01038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09588__A2 _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08154_ _03688_ _03689_ _03691_ _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__07599__A1 _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07105_ _02733_ _02736_ _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08085_ _03635_ _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07036_ _02614_ _02630_ _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05297_ _00970_ _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05058__I _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08987_ _04146_ _00594_ _04339_ _04343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07938_ ci_neuron.uut_simple_neuron.titan_id_2\[19\] ci_neuron.uut_simple_neuron.titan_id_5\[19\]
+ _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_3_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07869_ _03429_ _03432_ _03454_ _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_97_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09608_ _04789_ _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_39_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09539_ ci_neuron.output_val_internal\[24\] _04749_ _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09418__I3 _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09579__A2 _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_72_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09200__A1 _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08003__A2 ci_neuron.uut_simple_neuron.titan_id_5\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10245_ _00142_ net98 ci_neuron.uut_simple_neuron.titan_id_6\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10176_ _00073_ net211 ci_neuron.uut_simple_neuron.titan_id_2\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout190 net199 net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09503__A2 _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08562__I0 _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05220_ _00740_ _00896_ _00897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05151_ _00806_ _00827_ _00829_ _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06253__A1 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05082_ _00733_ _00753_ _00757_ _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_85_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08910_ internal_ih.byte4\[0\] internal_ih.byte3\[0\] _04296_ _04299_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09890_ _00051_ net23 ci_neuron.value_i\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08841_ internal_ih.byte0\[2\] _04254_ _04260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05984_ _01550_ _01641_ _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08772_ _03979_ _04218_ _04219_ _00303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07505__A1 _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07723_ ci_neuron.uut_simple_neuron.titan_id_4\[14\] ci_neuron.uut_simple_neuron.titan_id_3\[14\]
+ _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04935_ _00639_ _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07654_ ci_neuron.uut_simple_neuron.titan_id_4\[2\] ci_neuron.uut_simple_neuron.titan_id_3\[2\]
+ _03277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06605_ _02245_ _02202_ _02246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04866_ internal_ih.byte4\[3\] internal_ih.byte3\[3\] _00608_ _00614_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_36_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07585_ _03155_ _03210_ _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06536_ _02138_ _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09324_ _04574_ _00500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06467_ _01985_ _02109_ _02110_ _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09255_ _04531_ _00474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05418_ _00940_ _01011_ _01007_ _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_62_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08206_ net37 ci_neuron.uut_simple_neuron.x0\[1\] ci_neuron.uut_simple_neuron.x0\[2\]
+ _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06398_ _02006_ _02010_ _02042_ _02043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09186_ _03947_ _04489_ _04492_ _00444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07268__I _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05349_ _01010_ _01021_ _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08137_ ci_neuron.uut_simple_neuron.titan_id_1\[22\] ci_neuron.uut_simple_neuron.titan_id_0\[22\]
+ _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06244__A1 _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06172__I ci_neuron.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08068_ ci_neuron.uut_simple_neuron.titan_id_1\[10\] ci_neuron.uut_simple_neuron.titan_id_0\[10\]
+ _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07019_ _02593_ _02650_ _02651_ _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10030_ _00515_ net133 internal_ih.data_pointer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10228_ _00155_ net196 ci_neuron.uut_simple_neuron.titan_id_6\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10159_ ci_neuron.uut_simple_neuron.titan_id_0\[1\] net187 ci_neuron.uut_simple_neuron.titan_id_2\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08535__I0 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08160__A1 _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07370_ _02950_ _02960_ _02997_ _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_33_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06321_ _01896_ _01967_ _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_127_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06252_ _01873_ _01900_ _01901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09040_ _04385_ _04386_ _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05203_ _00751_ _00842_ _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06183_ _01834_ _01835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_96_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06226__A1 _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05134_ _00813_ _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05065_ _00748_ _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09942_ _00457_ net176 ci_neuron.uut_simple_neuron.x0\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09873_ _00064_ net30 ci_neuron.value_i\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08824_ _01754_ _04236_ _04249_ _00325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08755_ _04207_ _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07706_ _03319_ _03320_ _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05967_ _01611_ _01625_ _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05898_ _01557_ _01541_ _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08686_ _04152_ _04149_ _04153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04918_ _00648_ _00004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__04960__A1 internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07637_ _03197_ _03208_ _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04849_ _00594_ _00599_ _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07568_ _03157_ _03193_ _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06519_ _02158_ _02161_ _02162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09307_ _04564_ _00493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07499_ _03124_ _03125_ _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_11_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08454__A2 _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09238_ _04079_ _04503_ _04522_ _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09169_ ci_neuron.uut_simple_neuron.titan_id_6\[28\] _04481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10013_ ci_neuron.input_memory\[1\]\[13\] net173 ci_neuron.uut_simple_neuron.titan_id_1\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04951__A1 internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08445__A2 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_78_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07956__A1 _03512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ _02188_ _02337_ _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_05821_ _01368_ _01381_ _01480_ _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05752_ _01412_ _01391_ _01414_ _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_82_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08540_ _03968_ _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05683_ _01218_ _01325_ _01347_ _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_77_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08471_ _03968_ _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_46_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07422_ _03047_ _03049_ _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07353_ _02913_ _02982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07284_ _02846_ _02913_ _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06304_ _01949_ _01937_ _01950_ _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06235_ _01827_ _01884_ _01885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09023_ _04356_ _04364_ _04369_ _04370_ _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_115_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06166_ _01819_ _01820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05117_ _00734_ _00792_ _00797_ _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_06097_ _01750_ _01752_ _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05048_ net38 _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09925_ _00030_ net10 ci_neuron.instruction_i\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09856_ _00435_ net102 ci_neuron.output_memory\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07175__A2 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05066__I _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08807_ _04240_ _00317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06999_ _02606_ _02632_ _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09787_ _00366_ net56 internal_ih.byte4\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08738_ internal_ih.received_byte_count\[2\] _04195_ _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08669_ _04136_ _04137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06686__A1 _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08427__A2 _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09001__I net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06677__A1 _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08910__I0 internal_ih.byte4\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08418__A2 ci_neuron.uut_simple_neuron.x0\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06020_ _01568_ _01677_ _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07971_ ci_neuron.uut_simple_neuron.titan_id_2\[23\] ci_neuron.uut_simple_neuron.titan_id_5\[23\]
+ _03530_ _03538_ _03540_ _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_06922_ _02498_ _02556_ _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09710_ _00289_ net123 internal_ih.spi_rx_byte_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_06853_ _02181_ _02453_ _02488_ _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09641_ ci_neuron.stream_o\[22\] ci_neuron.output_memory\[22\] _04816_ _04819_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06784_ _02420_ _02368_ _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05804_ _01462_ _01463_ _01465_ _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_78_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09572_ ci_neuron.output_memory\[30\] _04766_ _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05735_ _01397_ _01398_ _01399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08523_ _04000_ _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08901__I0 internal_ih.byte3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05666_ _01292_ _01293_ _01330_ _01268_ _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_37_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07969__C ci_neuron.uut_simple_neuron.titan_id_5\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08454_ ci_neuron.value_i\[1\] _03953_ _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07405_ _02382_ _02947_ _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05597_ ci_neuron.uut_simple_neuron.x2\[19\] _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08385_ ci_neuron.uut_simple_neuron.x0\[27\] _03891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07336_ _02888_ _02894_ _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07267_ _02852_ _02896_ _02897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09006_ _04182_ _04354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07198_ _01907_ _02828_ _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06840__A1 _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06218_ _01860_ _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06149_ _01743_ _01796_ _01803_ _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09941__CLK net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09908_ _00004_ net7 ci_neuron.address_i\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09839_ _00418_ net195 ci_neuron.output_memory\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05331__A1 _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09620__I1 ci_neuron.output_memory\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05520_ _01147_ _01151_ _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05451_ _01121_ _00206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_117_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08170_ _03704_ _03705_ _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07075__A1 _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07121_ _02184_ _02691_ _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05382_ ci_neuron.uut_simple_neuron.x2\[12\] ci_neuron.uut_simple_neuron.x2\[13\]
+ ci_neuron.uut_simple_neuron.x2\[14\] _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_15_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07052_ _02339_ _02500_ _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_113_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06003_ _01462_ _01660_ _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09611__I1 ci_neuron.output_memory\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06050__A2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07954_ _03518_ _03523_ _03526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06905_ _02491_ _02510_ _02539_ _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07885_ _03462_ _03465_ _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06836_ _02470_ _02471_ _02472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09624_ ci_neuron.stream_o\[15\] ci_neuron.output_memory\[15\] _04805_ _04809_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06767_ _02401_ _02404_ _02405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_26_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09555_ _04746_ _04762_ _04763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06698_ _02228_ _02334_ _02336_ _02337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_78_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05718_ _01342_ _01381_ _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_53_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08506_ _03997_ _03998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09486_ _04704_ _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05649_ _01304_ _01314_ _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08437_ _03933_ _03937_ _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08368_ _03874_ _03875_ _03876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07319_ _02382_ _02947_ _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08299_ _03804_ _03805_ _03815_ _03803_ _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_18_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10261_ _00554_ net151 ci_neuron.stream_o\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08566__A1 _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09602__I1 ci_neuron.output_memory\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10192_ _00107_ net187 ci_neuron.uut_simple_neuron.titan_id_5\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07541__A2 ci_neuron.uut_simple_neuron.x3\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08766__S _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05552__A1 _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04951_ internal_ih.byte0\[2\] _00665_ _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_88_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07670_ ci_neuron.uut_simple_neuron.titan_id_4\[5\] ci_neuron.uut_simple_neuron.titan_id_3\[5\]
+ _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04882_ _00605_ _00625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06621_ _02215_ _02240_ _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05543__A1 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06552_ _02193_ _02194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09340_ _04566_ _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05503_ _01144_ _01154_ _01171_ _01132_ _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__09285__A2 _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09271_ _03933_ _04485_ _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_47_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06483_ _02100_ _02101_ _02126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08222_ _03729_ ci_neuron.uut_simple_neuron.x0\[5\] ci_neuron.uut_simple_neuron.x0\[4\]
+ _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05434_ _01104_ _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07048__A1 ci_neuron.uut_simple_neuron.x3\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05365_ _01036_ _01021_ _01037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08153_ ci_neuron.uut_simple_neuron.titan_id_1\[25\] ci_neuron.uut_simple_neuron.titan_id_0\[25\]
+ _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07104_ _02734_ _02735_ _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08084_ ci_neuron.uut_simple_neuron.titan_id_1\[13\] ci_neuron.uut_simple_neuron.titan_id_0\[13\]
+ _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07035_ _02661_ _02667_ _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05296_ _00969_ _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08986_ _00598_ _04340_ _04342_ _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07937_ _03508_ _03509_ _03511_ _03512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_48_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07868_ ci_neuron.uut_simple_neuron.titan_id_2\[3\] ci_neuron.uut_simple_neuron.titan_id_5\[3\]
+ _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07799_ _03396_ _03397_ _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06819_ _02452_ _02455_ _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09607_ _04799_ _00558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_39_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09538_ _04704_ _04749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09276__A2 _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09469_ _04673_ _04686_ _04688_ _04689_ _00530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_47_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10244_ _00141_ net98 ci_neuron.uut_simple_neuron.titan_id_6\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07211__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10175_ _00072_ net207 ci_neuron.uut_simple_neuron.titan_id_2\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout180 net181 net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout191 net194 net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08562__I1 _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07278__A1 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05150_ _00802_ _00825_ _00824_ _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05081_ _00735_ _00761_ _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09578__I0 ci_neuron.uut_simple_neuron.x0\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08840_ _04259_ _00331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05983_ _01597_ _01637_ _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08771_ _00795_ _04214_ _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07722_ _03330_ _03332_ _03333_ _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_04934_ _00657_ _00011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07653_ _03276_ _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04865_ _00613_ _00027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06604_ _02199_ _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07584_ _03194_ _03209_ _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09323_ _04069_ ci_neuron.input_memory\[1\]\[20\] _04572_ _04574_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07269__A1 _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06535_ _01856_ _02176_ _02177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06466_ _02036_ _02061_ _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09254_ _04119_ _03916_ _04490_ _04531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05417_ _01083_ _01086_ _01087_ _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08205_ _03729_ _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09185_ _03725_ _04491_ _04492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06397_ _02040_ _02041_ _02042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08769__A1 _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08136_ _03677_ _00078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05348_ _01012_ _01000_ _01020_ _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_114_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06244__A2 _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05279_ _00952_ _00953_ _00954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_70_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08067_ _03620_ _00094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07018_ _02596_ _02633_ _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08969_ _04192_ _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10227_ _00154_ net195 ci_neuron.uut_simple_neuron.titan_id_6\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10158_ ci_neuron.uut_simple_neuron.titan_id_0\[0\] net185 ci_neuron.uut_simple_neuron.titan_id_2\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10089_ _00186_ net77 ci_neuron.uut_simple_neuron.titan_id_0\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08535__I1 _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07922__I _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06320_ _01963_ _01966_ _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_57_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06251_ _01878_ _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05202_ _00855_ _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06182_ ci_neuron.uut_simple_neuron.x3\[0\] _01822_ _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_96_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07423__A1 _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05133_ _00812_ _00813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05064_ _00747_ _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_13_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09941_ _00456_ net172 ci_neuron.uut_simple_neuron.x0\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout83_I net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09872_ _00063_ net33 ci_neuron.value_i\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08823_ _04104_ _04237_ _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05966_ _01616_ _01624_ _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08754_ _03937_ _04206_ _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07705_ ci_neuron.uut_simple_neuron.titan_id_4\[10\] ci_neuron.uut_simple_neuron.titan_id_3\[10\]
+ ci_neuron.uut_simple_neuron.titan_id_4\[9\] ci_neuron.uut_simple_neuron.titan_id_3\[9\]
+ _03320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_04917_ internal_ih.byte5\[4\] _00646_ _00647_ internal_ih.byte1\[4\] _00648_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05897_ _01252_ _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08685_ internal_ih.spi_rx_byte_i\[2\] _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07636_ _03200_ _03207_ _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04848_ _00598_ internal_ih.current_instruction\[3\] internal_ih.current_instruction\[2\]
+ _00592_ _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_07567_ _03181_ _03192_ _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06518_ _02073_ _02159_ _02160_ _02161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09306_ _04027_ ci_neuron.input_memory\[1\]\[13\] _04561_ _04564_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07498_ _01984_ _03048_ _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09237_ _03862_ _04496_ _04522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_11_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06449_ _01998_ _02050_ _02092_ _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06183__I _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09168_ _04480_ _00438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08119_ _03662_ _03663_ _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_56_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09099_ _04365_ _04440_ _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07965__A2 ci_neuron.uut_simple_neuron.titan_id_5\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10012_ ci_neuron.input_memory\[1\]\[12\] net174 ci_neuron.uut_simple_neuron.titan_id_1\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08838__I _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05262__I _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07405__A1 _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05820_ _01477_ _01481_ _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_19_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05751_ _01413_ _01390_ _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05682_ _01331_ _01341_ _01346_ _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08470_ _03938_ _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07421_ _01984_ _03048_ _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_106_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_46_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07352_ _02846_ _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_92_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06303_ _01928_ _01948_ _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07283_ _02910_ _02912_ _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06234_ _01871_ _01883_ _01884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_86_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09022_ _04182_ _04370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_28_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06165_ ci_neuron.uut_simple_neuron.x3\[0\] _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05116_ _00794_ _00796_ _00797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07947__A2 ci_neuron.uut_simple_neuron.titan_id_5\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06096_ _00937_ _01751_ _01669_ _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09924_ _00029_ net9 ci_neuron.instruction_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05047_ _00715_ _00725_ _00732_ _00000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09855_ _00434_ net102 ci_neuron.output_memory\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08806_ _04064_ _01264_ _04239_ _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_0_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_37_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06998_ _02608_ _02631_ _02632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_99_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09786_ _00365_ net54 internal_ih.byte4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05949_ _01576_ _01585_ _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08737_ internal_ih.received_byte_count\[2\] _04195_ _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08668_ _04135_ _04136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07619_ _03181_ _03192_ _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08599_ _04076_ _04077_ _03953_ _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_91_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09870__CLK net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_46_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_55_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09560__A1 ci_neuron.output_memory\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08910__I1 internal_ih.byte3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09399__I _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_64_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09379__A1 ci_neuron.output_memory\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07970_ _03539_ _03540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06921_ ci_neuron.uut_simple_neuron.x3\[19\] _02555_ _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09551__A1 ci_neuron.output_memory\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06852_ _02182_ _02329_ _02488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_93_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09640_ _04818_ _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06783_ _01920_ _01938_ _02420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05803_ _01464_ _01431_ _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_78_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09571_ _04765_ _04773_ _04775_ _04776_ _00545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05734_ _00932_ _01351_ _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08522_ _03986_ _04010_ _04012_ _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08453_ _03925_ _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07404_ _02392_ _02946_ _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05665_ _00936_ _01329_ _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05596_ _01099_ _01102_ _01187_ _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_58_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08384_ _03889_ _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07335_ _02891_ _02893_ _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07266_ _02885_ _02895_ _02896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06217_ _01823_ _01867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09005_ _04351_ _04353_ _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07197_ _02273_ _02291_ _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06148_ _01621_ _01802_ _01803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06079_ _01648_ _01725_ _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08593__A2 _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09907_ _00003_ net13 ci_neuron.address_i\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09838_ _00417_ net193 ci_neuron.output_memory\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09769_ _00348_ net64 internal_ih.byte2\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06108__A1 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09012__I internal_ih.data_pointer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07084__A2 _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_72_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_129_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout250_I net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05450_ _01118_ _01120_ _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05381_ _00970_ _01005_ _01052_ _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07120_ _02190_ _02690_ _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07051_ _02502_ _02683_ _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06281__I _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06002_ _01374_ _01659_ _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_81_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07953_ ci_neuron.uut_simple_neuron.titan_id_2\[21\] ci_neuron.uut_simple_neuron.titan_id_5\[21\]
+ _03525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06904_ _02493_ _02509_ _02539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07884_ ci_neuron.uut_simple_neuron.titan_id_2\[9\] ci_neuron.uut_simple_neuron.titan_id_5\[9\]
+ _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06835_ _02365_ _02430_ _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09623_ _04808_ _00565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_90_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06766_ _02266_ _02402_ _02403_ _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09554_ _03892_ ci_neuron.input_memory\[1\]\[27\] _01706_ _03084_ _04760_ _04761_
+ _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_26_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06697_ _02335_ _02333_ _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05717_ ci_neuron.uut_simple_neuron.x2\[22\] _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_66_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08505_ _03769_ _03771_ _03987_ _03997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09485_ _04596_ _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05648_ _01313_ _01314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_92_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08436_ _03934_ _03936_ _03937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_93_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08367_ ci_neuron.uut_simple_neuron.x0\[25\] _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07318_ _02392_ _02946_ _02947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05579_ _01246_ _00209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08298_ ci_neuron.uut_simple_neuron.x0\[14\] ci_neuron.uut_simple_neuron.x0\[15\]
+ _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07249_ _02857_ _02878_ _02879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10260_ _00553_ net149 ci_neuron.stream_o\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08810__I0 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10191_ _00096_ net185 ci_neuron.uut_simple_neuron.titan_id_5\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09515__A1 ci_neuron.output_memory\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09054__I0 ci_neuron.output_val_internal\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04950_ _00667_ _00044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_88_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06620_ _02215_ _02240_ _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04881_ _00624_ _00032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08756__I _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10003__D ci_neuron.input_memory\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06551_ _01954_ _02192_ _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06482_ _01846_ _02125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05502_ _01058_ _01152_ _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09270_ _04540_ _04535_ _04541_ _00479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05433_ _01103_ _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08221_ ci_neuron.uut_simple_neuron.x0\[4\] ci_neuron.uut_simple_neuron.x0\[5\] _03733_
+ _03737_ _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_7_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07048__A2 ci_neuron.uut_simple_neuron.x3\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05364_ _01010_ _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_31_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08152_ _03690_ _00081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07103_ _02730_ ci_neuron.uut_simple_neuron.x3\[23\] _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05295_ ci_neuron.uut_simple_neuron.x2\[12\] _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08083_ ci_neuron.uut_simple_neuron.titan_id_1\[12\] ci_neuron.uut_simple_neuron.titan_id_0\[12\]
+ _03631_ _03632_ _03634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_113_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07034_ _02664_ _02666_ _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06559__A1 _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08985_ _04143_ _04341_ _04342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07936_ ci_neuron.uut_simple_neuron.titan_id_2\[18\] ci_neuron.uut_simple_neuron.titan_id_5\[18\]
+ _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07867_ ci_neuron.uut_simple_neuron.titan_id_2\[7\] ci_neuron.uut_simple_neuron.titan_id_5\[7\]
+ _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07798_ ci_neuron.uut_simple_neuron.titan_id_4\[27\] ci_neuron.uut_simple_neuron.titan_id_3\[27\]
+ _03397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06818_ _02454_ _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09606_ ci_neuron.stream_o\[7\] ci_neuron.output_memory\[7\] _04795_ _04799_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_39_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06749_ ci_neuron.uut_simple_neuron.x3\[15\] _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09537_ _04746_ _04747_ _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09468_ ci_neuron.output_val_internal\[14\] _04680_ _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08419_ _03919_ _03920_ _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09399_ _04602_ _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10243_ _00140_ net102 ci_neuron.uut_simple_neuron.titan_id_6\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10174_ _00071_ net206 ci_neuron.uut_simple_neuron.titan_id_2\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout181 net182 net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout192 net194 net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout170 net171 net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05080_ _00758_ _00759_ _00762_ _00161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05213__A1 _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05982_ _01640_ _00218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08770_ _04208_ _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07721_ ci_neuron.uut_simple_neuron.titan_id_4\[13\] ci_neuron.uut_simple_neuron.titan_id_3\[13\]
+ _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04933_ internal_ih.byte6\[3\] _00652_ _00653_ internal_ih.byte2\[3\] _00657_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07652_ ci_neuron.uut_simple_neuron.titan_id_4\[2\] ci_neuron.uut_simple_neuron.titan_id_3\[2\]
+ _03275_ _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_04864_ internal_ih.byte7\[2\] _00606_ _00612_ _00610_ _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06603_ _02241_ _02243_ _02244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_07583_ _03197_ _03208_ _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_36_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06534_ _01862_ _02175_ _02176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09322_ _04573_ _00499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07269__A2 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08466__A1 _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06465_ _02036_ _02061_ _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09253_ _04530_ _00473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06396_ _02005_ _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05416_ _01084_ _01085_ _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08204_ ci_neuron.uut_simple_neuron.x0\[3\] ci_neuron.uut_simple_neuron.x0\[4\] _03733_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_16_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09184_ _04490_ _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05347_ _01018_ _01019_ _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_71_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08135_ ci_neuron.uut_simple_neuron.titan_id_1\[22\] ci_neuron.uut_simple_neuron.titan_id_0\[22\]
+ _03676_ _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_16_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05278_ _00931_ _00933_ _00950_ _00953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08066_ _03618_ _03619_ _03620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07017_ _02596_ _02633_ _02650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09194__A2 _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08968_ _04331_ _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07919_ _03493_ _03495_ _03496_ _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_08899_ internal_ih.byte3\[3\] internal_ih.byte2\[3\] _04291_ _04293_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08457__A1 _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10226_ _00153_ net194 ci_neuron.uut_simple_neuron.titan_id_6\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10157_ _00222_ net235 ci_neuron.uut_simple_neuron.titan_id_3\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10088_ _00185_ net82 ci_neuron.uut_simple_neuron.titan_id_0\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout163_I net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08448__A1 _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06250_ _01898_ _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09248__I0 _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05201_ _00851_ _00875_ _00877_ _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08970__S _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06181_ _01833_ _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_96_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05132_ _00811_ _00812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05063_ ci_neuron.uut_simple_neuron.x2\[1\] _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09940_ _00455_ net168 ci_neuron.uut_simple_neuron.x0\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09871_ _00062_ net34 ci_neuron.value_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08822_ _01619_ _04236_ _04248_ _00324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05965_ _01617_ _01623_ _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08753_ _03934_ _03931_ _03928_ _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07704_ ci_neuron.uut_simple_neuron.titan_id_4\[10\] ci_neuron.uut_simple_neuron.titan_id_3\[10\]
+ _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04916_ _00627_ _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05896_ _01518_ _01554_ _01555_ _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08684_ internal_ih.spi_tx_byte_o\[1\] _04137_ _04142_ _04146_ _04151_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07635_ _03242_ _03245_ _03259_ _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_105_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04847_ internal_ih.current_instruction\[0\] _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_119_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07566_ _03184_ _03191_ _03192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06517_ _02108_ _02111_ _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09305_ _04563_ _00492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07497_ _02040_ _02009_ _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09236_ _04521_ _00465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06448_ _02089_ _02091_ _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_90_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06379_ _01981_ _02024_ _02023_ _02025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09167_ ci_neuron.uut_simple_neuron.titan_id_6\[27\] _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08118_ ci_neuron.uut_simple_neuron.titan_id_1\[19\] ci_neuron.uut_simple_neuron.titan_id_0\[19\]
+ _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_56_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09098_ ci_neuron.output_val_internal\[30\] ci_neuron.output_val_internal\[22\] ci_neuron.output_val_internal\[14\]
+ ci_neuron.output_val_internal\[6\] _04366_ _04367_ _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08049_ ci_neuron.uut_simple_neuron.titan_id_1\[7\] ci_neuron.uut_simple_neuron.titan_id_0\[7\]
+ _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_116_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10011_ ci_neuron.input_memory\[1\]\[11\] net253 ci_neuron.uut_simple_neuron.titan_id_1\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06925__A1 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_129_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08602__A1 _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07169__A1 ci_neuron.uut_simple_neuron.x3\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10209_ _00105_ net230 ci_neuron.uut_simple_neuron.titan_id_5\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05750_ _01208_ _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05681_ _01330_ _01343_ _01345_ _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07420_ _01997_ _02008_ _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_46_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07351_ _02840_ _02914_ _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06302_ _01928_ _01948_ _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07282_ _02781_ _02834_ _02911_ _02912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08841__A1 internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06233_ _01882_ _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_100_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09021_ _04365_ _04368_ _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06164_ _01818_ _00222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05115_ _00756_ _00766_ _00795_ _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06095_ ci_neuron.uut_simple_neuron.x2\[29\] _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09923_ _00028_ net10 ci_neuron.instruction_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05046_ _00715_ _00731_ ci_neuron.stream_enabled _00732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09854_ _00433_ net102 ci_neuron.output_memory\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08805_ _04224_ _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06997_ _02612_ _02614_ _02630_ _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09785_ _00364_ net56 internal_ih.byte4\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05948_ _01605_ _01606_ _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08736_ _04190_ _04194_ _04195_ _00291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05879_ _01464_ _01483_ _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08667_ spi_interface_cvonk.SCLK_r\[2\] _04125_ _04128_ _04135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_07618_ _03159_ _03180_ _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07883__A2 ci_neuron.uut_simple_neuron.titan_id_5\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08598_ _03861_ _04072_ _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07549_ _03162_ _03174_ _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_101_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09219_ _04034_ _03809_ _04509_ _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08435__I1 _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08849__I _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_110_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05885__A1 _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07874__A2 ci_neuron.uut_simple_neuron.titan_id_5\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08823__A1 _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09466__I3 _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05637__A1 _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07928__I _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07149__B _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06920_ ci_neuron.uut_simple_neuron.x3\[20\] _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06851_ _02438_ _02485_ _02486_ _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07562__A1 _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06782_ _02364_ _02367_ _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05802_ _01428_ _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09570_ ci_neuron.output_val_internal\[29\] _04771_ _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05733_ _01319_ _01350_ _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08521_ _02091_ _04011_ _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08452_ _03951_ _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_07403_ _03029_ _03030_ _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_102_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05664_ _01328_ _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05595_ _01192_ _01224_ _01228_ _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08383_ ci_neuron.uut_simple_neuron.x0\[26\] _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07334_ _01895_ _02313_ _02905_ _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_45_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07265_ _02888_ _02894_ _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_116_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06216_ _01866_ _00165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09004_ _04352_ _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07196_ _02825_ _02746_ _02826_ _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06147_ _01798_ _01801_ _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_113_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06078_ _01691_ _01724_ _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09906_ _00002_ net13 ci_neuron.address_i\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05029_ _00710_ _00714_ _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07553__A1 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09837_ _00416_ net193 ci_neuron.output_memory\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09768_ _00347_ net65 internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08719_ _04177_ _04179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_29_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09699_ spi_interface_cvonk.SS_r\[0\] net120 spi_interface_cvonk.SS_r\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_124_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07856__A2 ci_neuron.uut_simple_neuron.titan_id_5\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10075__CLK net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_75_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05380_ ci_neuron.uut_simple_neuron.x2\[14\] _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07050_ _02680_ _02682_ _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06283__A1 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06001_ _01614_ _01615_ _01658_ _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_70_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07607__B ci_neuron.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07952_ _03524_ _00140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06903_ _02531_ _02537_ _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07883_ ci_neuron.uut_simple_neuron.titan_id_2\[8\] ci_neuron.uut_simple_neuron.titan_id_5\[8\]
+ _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06834_ _02425_ _02426_ _02429_ _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08583__I0 _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ ci_neuron.stream_o\[14\] ci_neuron.output_memory\[14\] _04805_ _04808_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09553_ _03935_ _04761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06765_ _02311_ _02349_ _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_26_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08504_ _03951_ _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06696_ _02283_ _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05716_ _01379_ _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09484_ _04701_ _04702_ _04703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05647_ _01306_ _01307_ _01312_ _01313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_19_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08435_ ci_neuron.normalised_stream_write_address\[1\] _03935_ _03927_ _03936_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08366_ ci_neuron.uut_simple_neuron.x0\[24\] _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07317_ _02547_ _02876_ _02875_ _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05578_ _01240_ _01245_ _01246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07996__C ci_neuron.uut_simple_neuron.titan_id_5\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08297_ ci_neuron.uut_simple_neuron.x0\[15\] ci_neuron.uut_simple_neuron.x0\[16\]
+ _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__09460__A1 ci_neuron.output_memory\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07248_ _02873_ _02877_ _02878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07179_ _02617_ _02737_ _02809_ _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09212__A1 _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10190_ ci_neuron.uut_simple_neuron.titan_id_3\[0\] net183 ci_neuron.uut_simple_neuron.titan_id_5\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06577__A2 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08810__I1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07526__A1 _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09279__A1 _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05068__A2 _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04880_ internal_ih.byte7\[7\] _00616_ _00623_ _00597_ _00624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06550_ _01933_ _02049_ _02192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_48_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06481_ _02080_ _02106_ _02123_ _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_87_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05501_ _01137_ _01143_ _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05432_ _01099_ _01102_ _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08220_ ci_neuron.uut_simple_neuron.x0\[5\] ci_neuron.uut_simple_neuron.x0\[6\] _03747_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_56_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05363_ _00743_ _01008_ _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_31_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08151_ _03688_ _03689_ _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_125_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07102_ _02623_ _02734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05294_ _00863_ _00967_ _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08082_ _03633_ _00067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07033_ _01862_ _02665_ _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06559__A2 _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08984_ _04339_ _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07935_ _03510_ _00136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09605_ _04798_ _00557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07866_ _03452_ _00156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07797_ ci_neuron.uut_simple_neuron.titan_id_4\[26\] ci_neuron.uut_simple_neuron.titan_id_3\[26\]
+ _03395_ _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06817_ _02181_ _02453_ _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06748_ _02335_ _02338_ _02385_ _02386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_78_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09536_ _03877_ ci_neuron.input_memory\[1\]\[24\] _01475_ _02865_ _04738_ _04739_
+ _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_109_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09467_ _04677_ _04687_ _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06679_ _02316_ _02317_ _02318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08418_ ci_neuron.uut_simple_neuron.x0\[30\] ci_neuron.uut_simple_neuron.x0\[31\]
+ _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09398_ ci_neuron.output_memory\[4\] _04628_ _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08349_ _03856_ _03859_ _03860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_129_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05470__A2 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10242_ _00139_ net104 ci_neuron.uut_simple_neuron.titan_id_6\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08795__I0 _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10173_ _00070_ net267 ci_neuron.uut_simple_neuron.titan_id_2\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09018__I internal_ih.data_pointer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout182 net215 net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout160 net161 net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout171 net172 net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout193 net194 net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09424__A1 ci_neuron.output_memory\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09578__I2 ci_neuron.uut_simple_neuron.x2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08786__I0 _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05981_ _01637_ _01639_ _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07720_ ci_neuron.uut_simple_neuron.titan_id_4\[13\] ci_neuron.uut_simple_neuron.titan_id_3\[13\]
+ _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_04932_ _00656_ _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07651_ ci_neuron.uut_simple_neuron.titan_id_4\[1\] ci_neuron.uut_simple_neuron.titan_id_3\[1\]
+ _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04863_ internal_ih.byte4\[2\] internal_ih.byte3\[2\] _00608_ _00612_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07582_ _03200_ _03207_ _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06602_ _02170_ _02198_ _02242_ _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_88_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06533_ _01926_ _02044_ _02174_ _02175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09321_ _04064_ ci_neuron.input_memory\[1\]\[19\] _04572_ _04573_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_36_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06464_ _02075_ _02077_ _02107_ _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_90_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09252_ _04116_ _03915_ _04490_ _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06395_ _01997_ _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05415_ _01084_ _01085_ _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_16_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09415__A1 ci_neuron.output_memory\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09183_ _04487_ _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08203_ _03732_ _00193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05346_ _01002_ _00983_ _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_71_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08134_ _03672_ _03673_ _03675_ _03676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_43_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05277_ _00951_ _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08065_ ci_neuron.uut_simple_neuron.titan_id_1\[10\] ci_neuron.uut_simple_neuron.titan_id_0\[10\]
+ _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07016_ _01831_ _02592_ _02649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08967_ internal_ih.byte7\[1\] internal_ih.byte6\[1\] _04327_ _04331_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07918_ ci_neuron.uut_simple_neuron.titan_id_2\[15\] ci_neuron.uut_simple_neuron.titan_id_5\[15\]
+ _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08898_ _04292_ _00356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07849_ _03434_ _03435_ _03438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09519_ _04721_ _04729_ _04731_ _04732_ _00537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__08457__A2 _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10225_ _00152_ net159 ci_neuron.uut_simple_neuron.titan_id_6\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10156_ _00221_ net235 ci_neuron.uut_simple_neuron.titan_id_3\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10087_ _00184_ net82 ci_neuron.uut_simple_neuron.titan_id_0\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout156_I net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05200_ _00854_ _00874_ _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06180_ _01832_ _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_96_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05131_ ci_neuron.uut_simple_neuron.x2\[6\] _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05062_ _00746_ _00159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09870_ _00061_ net34 ci_neuron.value_i\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08821_ _04099_ _04237_ _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05964_ _01621_ _01622_ _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08752_ _04194_ _04205_ _00297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout69_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07703_ _03313_ _03316_ _03318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08683_ _04134_ _04144_ _04150_ _00283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04915_ _00639_ _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07634_ _03010_ _03248_ _03258_ _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__06698__A1 _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05895_ _01520_ _01543_ _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04846_ _00596_ _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07565_ _03190_ _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07496_ _03121_ _03122_ _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06516_ _02108_ _02111_ _02159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_91_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09304_ _04023_ ci_neuron.input_memory\[1\]\[12\] _04561_ _04563_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06447_ _02090_ _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09235_ _04074_ _03851_ _04519_ _04521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_106_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06378_ _01943_ _01979_ _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09166_ _04479_ _00437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05329_ _00970_ _00940_ _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08117_ _03660_ _03661_ _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09097_ _04417_ ci_neuron.stream_o\[6\] ci_neuron.stream_o\[22\] _04418_ _04438_
+ _04439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XTAP_TAPCELL_ROW_56_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08048_ ci_neuron.uut_simple_neuron.titan_id_1\[7\] ci_neuron.uut_simple_neuron.titan_id_0\[7\]
+ ci_neuron.uut_simple_neuron.titan_id_1\[6\] ci_neuron.uut_simple_neuron.titan_id_0\[6\]
+ _03604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_31_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07178__A2 _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10010_ ci_neuron.input_memory\[1\]\[10\] net255 ci_neuron.uut_simple_neuron.titan_id_1\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09999_ _00514_ net129 internal_ih.expected_byte_count\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06925__A2 _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_67_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08602__A2 _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09650__I1 ci_neuron.output_memory\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07169__A2 ci_neuron.uut_simple_neuron.x3\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10208_ _00104_ net282 ci_neuron.uut_simple_neuron.titan_id_5\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10139_ _00204_ net277 ci_neuron.uut_simple_neuron.titan_id_3\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04927__B2 internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05680_ _00740_ _01344_ _01329_ _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07350_ _02916_ _02978_ _02979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06301_ _01935_ _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07281_ _02784_ _02833_ _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05104__A1 _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08841__A2 _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09020_ ci_neuron.output_val_internal\[24\] ci_neuron.output_val_internal\[16\] ci_neuron.output_val_internal\[8\]
+ ci_neuron.output_val_internal\[0\] _04366_ _04367_ _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_115_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06232_ _01829_ _01881_ _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_100_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08780__I _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06163_ _01807_ _01815_ _01817_ _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09967__CLK net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05114_ _00793_ _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09641__I1 ci_neuron.output_memory\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06094_ _01714_ _01715_ _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09922_ _00027_ net10 ci_neuron.instruction_i\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_05045_ _00728_ _00730_ _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09853_ _00432_ net103 ci_neuron.output_memory\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08804_ _01266_ _04236_ _04238_ _00316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09784_ _00363_ net48 internal_ih.byte4\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06996_ _02619_ _02627_ _02629_ _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_56_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08735_ internal_ih.received_byte_count\[1\] _04189_ _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05947_ _01567_ _01588_ _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05878_ _01464_ _01483_ _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08666_ _04133_ _04134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07617_ _03240_ _03241_ _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08597_ _03862_ _04072_ _04076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07548_ _03172_ _03173_ _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07479_ _03105_ _03106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_62_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09218_ _04511_ _00457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09149_ ci_neuron.uut_simple_neuron.titan_id_6\[18\] _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09632__I1 ci_neuron.output_memory\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04909__A1 internal_ih.byte5\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04909__B2 internal_ih.byte1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08823__A2 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08533__C _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout119_I net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06850_ _02440_ _02456_ _02486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05801_ _01428_ _01431_ _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08976__S _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06781_ _02359_ _02416_ _02417_ _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05732_ _00932_ _01395_ _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08775__I _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08520_ _03939_ _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10022__D ci_neuron.input_memory\[1\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05663_ _01327_ _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08511__A1 _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08451_ _03950_ _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07402_ _01969_ _02957_ _03030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_102_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05594_ _01083_ _01210_ _01176_ _01260_ _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08382_ _03888_ _00186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07333_ _02922_ _02961_ _02962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_116_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07264_ _02891_ _02893_ _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_60_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06215_ _01851_ _01865_ _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09003_ _04173_ _04174_ _04181_ _04192_ _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_26_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07195_ _02276_ _02745_ _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06146_ _01699_ _01799_ _01800_ _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_113_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06077_ _01733_ _00220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09905_ _00024_ net14 ci_neuron.address_i\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05028_ ci_neuron.instruction_i\[0\] ci_neuron.instruction_i\[1\] _00713_ _00714_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09836_ _00415_ net191 ci_neuron.output_memory\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06979_ _02550_ _02559_ _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09767_ _00346_ net65 internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08718_ internal_ih.instruction_received _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09698_ net2 net120 spi_interface_cvonk.SS_r\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08502__A1 _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08649_ _04119_ ci_neuron.uut_simple_neuron.x3\[30\] _04111_ _04120_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_64_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09302__I0 _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07480__A1 _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06000_ _01580_ _01613_ _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07951_ _03522_ _03523_ _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06902_ _02534_ _02536_ _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07882_ _03466_ _00158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06833_ _02469_ _00237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08583__I1 _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09621_ _04807_ _00564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06764_ _02311_ _02349_ _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_78_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09552_ _03930_ _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_fanout51_I net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05715_ ci_neuron.uut_simple_neuron.x2\[21\] ci_neuron.uut_simple_neuron.x2\[22\]
+ _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08503_ _03986_ _03994_ _03995_ _00258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09288__A2 _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06695_ _02283_ _02333_ _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09483_ _03822_ ci_neuron.input_memory\[1\]\[16\] _01150_ _02384_ _04691_ _04692_
+ _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_59_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05646_ _01309_ _01277_ _01311_ _01312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_92_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08434_ ci_neuron.address_i\[1\] _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05577_ _01243_ _01244_ _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08365_ _03873_ _00184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07316_ _02926_ _02944_ _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08296_ _03813_ _00175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06274__A2 _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07247_ _02547_ _02876_ _02877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07178_ _02808_ _02736_ _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09212__A2 _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06129_ _01743_ _01775_ _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09819_ _00398_ net58 internal_ih.current_instruction\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_126_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07214__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09214__I _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06480_ _02084_ _02105_ _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05500_ _01130_ _01167_ _01168_ _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05431_ _01100_ _01101_ _00963_ _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_28_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08150_ ci_neuron.uut_simple_neuron.titan_id_1\[25\] ci_neuron.uut_simple_neuron.titan_id_0\[25\]
+ _03689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_07101_ _02620_ _02681_ _02732_ _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_99_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05362_ _00888_ _00985_ _01033_ _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_31_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05293_ _00891_ _00914_ _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08081_ _03631_ _03632_ _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_31_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07032_ _02175_ _02193_ _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08983_ _04339_ _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07934_ _03508_ _03509_ _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07865_ _03450_ _03451_ _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_3_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09604_ ci_neuron.stream_o\[6\] ci_neuron.output_memory\[6\] _04795_ _04798_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07796_ _03387_ _03388_ _03394_ _03391_ _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06816_ _02144_ _02285_ _02453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_78_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06747_ _02333_ _02384_ _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09535_ _04700_ _04746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_39_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06678_ _01891_ _01938_ _02317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09466_ _03809_ ci_neuron.input_memory\[1\]\[14\] _01052_ _02335_ _04667_ _04669_
+ _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_121_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05629_ _01288_ _01294_ _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08417_ _03917_ _03918_ _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_50_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09397_ _04599_ _04628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08348_ _03844_ _03846_ _03857_ _03858_ _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_46_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08279_ _03795_ _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05099__I _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10241_ _00137_ net69 ci_neuron.uut_simple_neuron.titan_id_6\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10172_ _00069_ net268 ci_neuron.uut_simple_neuron.titan_id_2\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout172 net182 net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout150 net163 net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout161 net162 net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout183 net185 net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout194 net198 net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09188__A1 _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout101_I net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05980_ _01597_ _01598_ _01638_ _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04931_ internal_ih.byte6\[2\] _00652_ _00653_ internal_ih.byte2\[2\] _00656_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07650_ _03274_ _00249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04862_ _00611_ _00026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07581_ _01833_ _03206_ _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06601_ _02172_ _02197_ _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06532_ _02173_ _02148_ _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09320_ _04566_ _04572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09502__I3 _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09251_ _04529_ _00472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06463_ _02080_ _02106_ _02107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08202_ _03726_ _03730_ _03731_ _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06394_ _01867_ _02038_ _02039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05414_ _01047_ _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09182_ _04488_ _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05345_ _01017_ _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08133_ ci_neuron.uut_simple_neuron.titan_id_1\[21\] ci_neuron.uut_simple_neuron.titan_id_0\[21\]
+ _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08064_ _03614_ _03616_ _03617_ _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_31_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07015_ _02639_ _02637_ _02647_ _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05276_ _00931_ _00933_ _00950_ _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08966_ _04330_ _00386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07917_ ci_neuron.uut_simple_neuron.titan_id_2\[15\] ci_neuron.uut_simple_neuron.titan_id_5\[15\]
+ _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08897_ internal_ih.byte3\[2\] internal_ih.byte2\[2\] _04291_ _04292_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07848_ ci_neuron.uut_simple_neuron.titan_id_2\[4\] ci_neuron.uut_simple_neuron.titan_id_5\[4\]
+ _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07779_ _03379_ _03380_ _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09518_ ci_neuron.output_val_internal\[21\] _04727_ _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09449_ _04649_ _04665_ _04671_ _04672_ _00527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_124_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10224_ _00149_ net191 ci_neuron.uut_simple_neuron.titan_id_6\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10155_ _00220_ net236 ci_neuron.uut_simple_neuron.titan_id_3\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08868__I _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10086_ _00183_ net95 ci_neuron.uut_simple_neuron.titan_id_0\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07408__A1 _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05130_ _00808_ _00809_ _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07959__A2 ci_neuron.uut_simple_neuron.titan_id_5\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08081__A1 _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04890__B2 internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05061_ _00737_ _00745_ _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08820_ _04247_ _00323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05963_ ci_neuron.uut_simple_neuron.x2\[1\] ci_neuron.uut_simple_neuron.x2\[27\]
+ _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08751_ internal_ih.received_byte_count\[7\] _04204_ _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05894_ _01520_ _01543_ _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07702_ _03317_ _00126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04914_ _00645_ _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08682_ _04146_ _04149_ _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07633_ _03251_ _03254_ _03257_ _03258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_04845_ internal_ih.current_instruction\[3\] _00592_ _00593_ _00595_ _00596_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07564_ _03187_ _03189_ _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_105_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07495_ _03031_ _03037_ _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06515_ _02154_ _02157_ _02158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09303_ _04562_ _00491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06446_ ci_neuron.uut_simple_neuron.x3\[10\] _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09234_ _04520_ _00464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09165_ ci_neuron.uut_simple_neuron.titan_id_6\[26\] _04479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06377_ _02016_ _02022_ _02023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08116_ _03657_ _03658_ _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05328_ _00892_ _01000_ _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_71_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09096_ _04405_ _04437_ _04438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05259_ _00905_ _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_56_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08047_ _03594_ _03599_ _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09411__I2 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__A1 _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09998_ _00513_ net129 internal_ih.expected_byte_count\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08949_ internal_ih.byte6\[1\] internal_ih.byte5\[1\] _04317_ _04321_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08637__B _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05287__I _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10207_ _00103_ net278 ci_neuron.uut_simple_neuron.titan_id_5\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10138_ _00203_ net277 ci_neuron.uut_simple_neuron.titan_id_3\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06129__A1 _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10069_ _00196_ net202 ci_neuron.uut_simple_neuron.titan_id_0\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout266_I net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05750__I _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07280_ _02847_ _02850_ _02909_ _02910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06300_ _01946_ _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06231_ _01877_ _01880_ _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_73_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06162_ _01779_ _01781_ _01816_ _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06093_ _01747_ _01748_ _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05113_ _00756_ _00766_ _00793_ _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_41_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09921_ _00026_ net24 ci_neuron.instruction_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05044_ _00708_ _00729_ _00713_ _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_111_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06368__A1 _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09852_ _00431_ net168 ci_neuron.output_memory\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08803_ _04059_ _04237_ _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09783_ _00362_ net47 internal_ih.byte4\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06995_ _02329_ _02628_ _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08734_ _04193_ _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05946_ _01572_ _01587_ _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05877_ _01523_ _01537_ _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08665_ _04124_ _04133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07616_ _02550_ _03178_ _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08596_ _04075_ _00271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07547_ _02733_ _02736_ _03012_ _03173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_48_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07478_ _03078_ _03104_ _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_62_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06429_ _02013_ _02031_ _02012_ _02062_ _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_63_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09217_ _04027_ _03797_ _04509_ _04511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09148_ _04470_ _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09079_ ci_neuron.output_val_internal\[28\] ci_neuron.output_val_internal\[20\] ci_neuron.output_val_internal\[12\]
+ ci_neuron.output_val_internal\[4\] _04390_ _04391_ _04423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__07020__A2 _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_129_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_24_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_33_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08587__A2 _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08831__I0 _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05270__A1 _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05800_ _01461_ _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_42_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06780_ _02361_ _02400_ _02417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05731_ _01359_ _01394_ _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05662_ _01326_ _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08450_ _03934_ _03950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07401_ _02374_ _02395_ _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_102_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08381_ _03886_ _03887_ _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07332_ _02950_ _02960_ _02961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05593_ _00887_ _01210_ _01211_ _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__07078__A2 _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07263_ _01935_ _02892_ _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_51_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07194_ _02225_ _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06214_ _01857_ _01864_ _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09002_ _04350_ _04254_ _04178_ _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06145_ _01746_ _01770_ _01699_ _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06589__A1 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06076_ _01729_ _01732_ _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05027_ ci_neuron.instruction_i\[2\] _00711_ _00712_ _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_09904_ _00023_ net13 ci_neuron.address_i\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_60_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09835_ _00414_ net160 ci_neuron.output_memory\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05013__A1 internal_ih.byte3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06978_ _02178_ _02611_ _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09766_ _00345_ net67 internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05929_ _01568_ _01588_ _01589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08717_ _04173_ _04176_ internal_ih.instruction_received _04177_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09697_ spi_interface_cvonk.SCLK_r\[1\] net120 spi_interface_cvonk.SCLK_r\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08648_ ci_neuron.value_i\[30\] _04118_ _04026_ _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08579_ _03840_ _04044_ _03852_ _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05004__A1 internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06752__A1 _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06396__I _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09500__I _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05491__A1 _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07950_ ci_neuron.uut_simple_neuron.titan_id_2\[21\] ci_neuron.uut_simple_neuron.titan_id_5\[21\]
+ _03523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06901_ _01832_ _02535_ _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07881_ _03464_ _03465_ _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_37_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06832_ _02466_ _02468_ _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09620_ ci_neuron.stream_o\[13\] ci_neuron.output_memory\[13\] _04805_ _04807_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06763_ _02359_ _02361_ _02400_ _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09551_ ci_neuron.output_memory\[27\] _04744_ _04759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05714_ _01146_ _01376_ _01377_ _01378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08502_ _01998_ _03980_ _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06694_ ci_neuron.uut_simple_neuron.x3\[15\] _02333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09482_ _04700_ _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05645_ _01279_ _01310_ _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08433_ _03929_ _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05576_ _01123_ _01162_ _01200_ _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_46_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08364_ _03869_ _03872_ _03873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07315_ _02942_ _02943_ _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08295_ _03809_ _03810_ _03812_ _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_116_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07246_ _02874_ _02875_ _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07177_ _02726_ _02806_ _02807_ _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_42_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06128_ _01771_ _01774_ _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06059_ _01714_ _01715_ _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_6_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09818_ _00397_ net61 internal_ih.current_instruction\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_126_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09749_ _00328_ net90 ci_neuron.uut_simple_neuron.x2\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08629__C _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09320__I _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05473__A1 _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout179_I net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08478__A1 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05430_ _00969_ _01005_ ci_neuron.uut_simple_neuron.x2\[14\] _01101_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_74_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05361_ _01012_ _01020_ _01033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_16_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07100_ _02623_ _02731_ _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_31_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05292_ _00941_ _00943_ _00965_ _00916_ _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_70_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08080_ ci_neuron.uut_simple_neuron.titan_id_1\[12\] ci_neuron.uut_simple_neuron.titan_id_0\[12\]
+ _03632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07031_ _02662_ _02611_ _02663_ _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05216__A1 ci_neuron.uut_simple_neuron.x2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08982_ _04183_ _04185_ _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07933_ ci_neuron.uut_simple_neuron.titan_id_2\[18\] ci_neuron.uut_simple_neuron.titan_id_5\[18\]
+ _03509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_48_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07864_ ci_neuron.uut_simple_neuron.titan_id_2\[7\] ci_neuron.uut_simple_neuron.titan_id_5\[7\]
+ _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_3_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06815_ _02444_ _02451_ _02452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09603_ _04797_ _00556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07795_ ci_neuron.uut_simple_neuron.titan_id_4\[26\] ci_neuron.uut_simple_neuron.titan_id_3\[26\]
+ _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06746_ _02383_ _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09534_ ci_neuron.output_memory\[24\] _04744_ _04745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06677_ _01891_ _01938_ _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_38_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09465_ ci_neuron.output_memory\[14\] _04675_ _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_121_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05628_ _01292_ _01293_ _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08416_ _03910_ _03913_ _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09396_ _04597_ _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05559_ _01226_ _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08347_ _03836_ _03850_ ci_neuron.uut_simple_neuron.x0\[20\] _03858_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08278_ _03795_ _03797_ _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08641__A1 _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07229_ _02801_ _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_59_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10240_ _00136_ net158 ci_neuron.uut_simple_neuron.titan_id_6\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10171_ _00068_ net268 ci_neuron.uut_simple_neuron.titan_id_2\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xfanout140 net146 net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout173 net175 net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout151 net157 net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout162 net163 net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout184 net185 net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout195 net198 net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07380__A1 ci_neuron.uut_simple_neuron.x3\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Left_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09188__A2 _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_94_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04930_ _00655_ _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_04861_ internal_ih.byte7\[1\] _00606_ _00609_ _00610_ _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06600_ _02213_ _02215_ _02240_ _02241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07580_ _03203_ _03205_ _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06531_ _01925_ _02173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_36_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07123__A1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09250_ _04110_ _03904_ _04525_ _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06462_ _02084_ _02105_ _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_91_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08201_ _03724_ _03727_ _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06393_ _01853_ _01925_ _02037_ _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05413_ _01044_ _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09181_ _04487_ _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05344_ _00976_ _01015_ _01016_ _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_71_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08132_ _03674_ _00076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05275_ _00934_ _00949_ _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08063_ ci_neuron.uut_simple_neuron.titan_id_1\[9\] ci_neuron.uut_simple_neuron.titan_id_0\[9\]
+ ci_neuron.uut_simple_neuron.titan_id_1\[8\] ci_neuron.uut_simple_neuron.titan_id_0\[8\]
+ _03617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_3_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07014_ _02634_ _02636_ _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_102_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08965_ internal_ih.byte7\[0\] internal_ih.byte6\[0\] _04327_ _04330_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07916_ _03494_ _00133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08896_ _04290_ _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07847_ _03436_ _00153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07778_ _03376_ _03377_ _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10221__D _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06729_ _02366_ _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09517_ _04724_ _04730_ _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09448_ ci_neuron.output_val_internal\[11\] _04655_ _04672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09379_ ci_neuron.output_memory\[1\] _04600_ _04613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10223_ _00138_ net186 ci_neuron.uut_simple_neuron.titan_id_6\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10154_ _00219_ net237 ci_neuron.uut_simple_neuron.titan_id_3\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10085_ _00182_ net107 ci_neuron.uut_simple_neuron.titan_id_0\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout211_I net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05060_ _00744_ _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06919__A1 _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05962_ _01618_ _01620_ _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08750_ internal_ih.received_byte_count\[6\] _04202_ _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05893_ _01553_ _00216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07701_ _03315_ _03316_ _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08681_ _04148_ _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04913_ internal_ih.byte5\[3\] _00640_ _00641_ internal_ih.byte1\[3\] _00645_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07632_ _03255_ _03256_ _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04844_ _00594_ internal_ih.current_instruction\[2\] _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07563_ _02132_ _03188_ _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_105_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09302_ _04017_ ci_neuron.input_memory\[1\]\[11\] _04561_ _04562_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07494_ _03034_ _03036_ _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06514_ _02075_ _02155_ _02156_ _02157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_48_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06445_ _02001_ _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09233_ _04069_ _03849_ _04519_ _04520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09164_ _04478_ _00436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06376_ _02017_ _02020_ _02021_ _02022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08115_ ci_neuron.uut_simple_neuron.titan_id_1\[18\] ci_neuron.uut_simple_neuron.titan_id_0\[18\]
+ _03660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05327_ _00886_ _00914_ _00984_ _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09095_ _04419_ ci_neuron.stream_o\[14\] _04437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05258_ _00932_ _00921_ _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08046_ _03588_ _03591_ _03601_ _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_31_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_79_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05189_ ci_neuron.uut_simple_neuron.x2\[8\] _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08969__I _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09411__I3 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07583__A1 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09997_ _00512_ net132 internal_ih.expected_byte_count\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08948_ _04320_ _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08879_ _04281_ _00348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_67_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_88_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05568__I _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_97_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_78_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05821__A1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10126__D net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10206_ _00102_ net270 ci_neuron.uut_simple_neuron.titan_id_5\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09563__A2 _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10137_ _00202_ net277 ci_neuron.uut_simple_neuron.titan_id_3\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10068_ _00195_ net201 ci_neuron.uut_simple_neuron.titan_id_0\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07326__A1 _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06230_ _01838_ _01879_ _01880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_100_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06161_ _01737_ _01778_ _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06092_ _01663_ _01717_ _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05112_ ci_neuron.uut_simple_neuron.x2\[5\] _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05812__A1 _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09920_ _00025_ net24 ci_neuron.instruction_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05043_ _00709_ _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09851_ _00430_ net68 ci_neuron.output_memory\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06994_ _02286_ _02447_ _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08802_ _04207_ _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09782_ _00361_ net47 internal_ih.byte3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05945_ _01602_ _01603_ _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08733_ _04191_ _04192_ _04187_ _04188_ _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_05876_ _01527_ _01536_ _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08664_ _04130_ _04132_ _00282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07615_ _02559_ _03177_ _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08595_ _04074_ _02804_ _04053_ _04075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07546_ _03165_ _03171_ _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07477_ _03100_ _03103_ _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09216_ _04510_ _00456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06428_ _02029_ _02071_ _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_62_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06359_ _01926_ _02004_ _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_16_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09147_ ci_neuron.uut_simple_neuron.titan_id_6\[17\] _04470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06056__A1 _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09078_ _04417_ ci_neuron.stream_o\[4\] ci_neuron.stream_o\[20\] _04418_ _04421_
+ _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_31_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08029_ _03584_ _03586_ _03587_ _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_31_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07556__A1 _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07859__A2 ci_neuron.uut_simple_neuron.titan_id_5\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08831__I1 ci_neuron.uut_simple_neuron.x2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08595__I0 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05730_ _01361_ _01366_ _01393_ _01394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_89_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05661_ _01266_ _01290_ _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07400_ _03001_ _03027_ _03028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_102_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08380_ ci_neuron.uut_simple_neuron.x0\[25\] ci_neuron.uut_simple_neuron.x0\[26\]
+ _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07331_ _02953_ _02959_ _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05592_ _01221_ _01230_ _01258_ _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07262_ _02323_ _02344_ _02892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07193_ _02822_ _02823_ _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06213_ _01863_ _01864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09001_ net31 _04350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06144_ _01746_ _01770_ _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_5_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06075_ _01730_ _01731_ _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_113_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09903_ _00022_ net14 ci_neuron.address_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05026_ ci_neuron.instruction_i\[4\] ci_neuron.instruction_i\[7\] ci_neuron.instruction_i\[6\]
+ _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_1_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09834_ _00413_ net159 ci_neuron.output_memory\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06210__A1 _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06977_ _02146_ _02610_ _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_09765_ _00344_ net65 internal_ih.byte1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05928_ _01572_ _01587_ _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08716_ _04174_ _04175_ _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09696_ spi_interface_cvonk.SCLK_r\[0\] net120 spi_interface_cvonk.SCLK_r\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08889__I1 internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05859_ _01467_ _01486_ _01519_ _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_83_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08647_ _03916_ _03910_ _04107_ _04118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_64_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08578_ _04060_ _00268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07529_ _03154_ _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_92_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_75_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08577__I0 _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09254__S _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06504__A2 _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06900_ _02079_ _02102_ _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_128_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07880_ ci_neuron.uut_simple_neuron.titan_id_2\[9\] ci_neuron.uut_simple_neuron.titan_id_5\[9\]
+ _03465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06831_ _02467_ _02406_ _02410_ _02414_ _02468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_06762_ _02369_ _02399_ _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09550_ _04743_ _04755_ _04757_ _04758_ _00542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_37_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05713_ _01375_ _01336_ _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09481_ _00728_ _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08501_ ci_neuron.value_i\[8\] _03944_ _03993_ _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06693_ _02182_ _02287_ _02331_ _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_08432_ _03928_ _03932_ _03933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08496__A2 _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05644_ _01247_ _01308_ _01277_ _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_59_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05575_ _01241_ _01242_ _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08363_ _03866_ _03870_ _03871_ _03865_ _03872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_116_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07314_ _02554_ _02557_ _02733_ _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_74_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08294_ _03803_ _03806_ _03811_ _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07245_ _02548_ _02680_ _02875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_33_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07176_ _02804_ _02805_ _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06127_ _01782_ _00221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06431__A1 _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06058_ ci_neuron.uut_simple_neuron.x2\[29\] _01670_ _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05009_ _00700_ _00052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_6_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09817_ _00396_ net59 internal_ih.current_instruction\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_126_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09748_ _00327_ net89 ci_neuron.uut_simple_neuron.x2\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09679_ _00266_ net233 ci_neuron.uut_simple_neuron.x3\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06498__A1 _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_25_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05170__A1 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09436__A1 ci_neuron.output_memory\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09924__CLK net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04984__A1 internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05360_ _01001_ _01030_ _01031_ _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05291_ _00739_ _00964_ _00965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07030_ _02146_ _02610_ _02663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08981_ _04338_ _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07932_ ci_neuron.uut_simple_neuron.titan_id_2\[17\] ci_neuron.uut_simple_neuron.titan_id_5\[17\]
+ _03497_ _03505_ _03507_ _03508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_07863_ ci_neuron.uut_simple_neuron.titan_id_2\[6\] ci_neuron.uut_simple_neuron.titan_id_5\[6\]
+ _03449_ _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_3_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06814_ _02330_ _02450_ _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09602_ ci_neuron.stream_o\[5\] ci_neuron.output_memory\[5\] _04795_ _04797_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07794_ _03393_ _00113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09533_ _04674_ _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06745_ ci_neuron.uut_simple_neuron.x3\[16\] _02383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06676_ _02312_ _02314_ _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09464_ _04673_ _04682_ _04684_ _04685_ _00529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_121_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05627_ _01263_ _01267_ _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09395_ _04598_ _04621_ _04625_ _04626_ _00519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_08415_ _03915_ _03916_ _03917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08346_ ci_neuron.uut_simple_neuron.x0\[20\] ci_neuron.uut_simple_neuron.x0\[21\]
+ _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_50_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05558_ ci_neuron.uut_simple_neuron.x2\[18\] _01226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05489_ _01081_ _01113_ _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08277_ _03796_ _03797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10219__D _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07228_ _02799_ _02858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07159_ _02720_ _02748_ _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06404__A1 _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10170_ _00067_ net267 ci_neuron.uut_simple_neuron.titan_id_2\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout130 net134 net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout174 net175 net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout152 net157 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout141 net145 net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout163 net164 net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout185 net190 net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout196 net197 net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07380__A2 ci_neuron.uut_simple_neuron.x3\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06955__I _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09331__I _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08632__A2 _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_108_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout289_I net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04860_ _00596_ _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06530_ _02134_ _02150_ _02171_ _02172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06461_ _02099_ _02104_ _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05412_ _00887_ _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08200_ _03729_ _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_117_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06392_ _01852_ _02007_ _02037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09180_ _04486_ _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05343_ _01013_ _01014_ _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08131_ _03672_ _03673_ _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08623__A2 _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06634__A1 _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05274_ _00935_ _00948_ _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08062_ _03606_ _03615_ _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07013_ _02646_ _00240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08964_ _04329_ _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_126_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07915_ ci_neuron.uut_simple_neuron.titan_id_2\[15\] ci_neuron.uut_simple_neuron.titan_id_5\[15\]
+ _03493_ _03494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09416__I _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08895_ _04256_ _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07846_ _03434_ _03435_ _03436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07777_ ci_neuron.uut_simple_neuron.titan_id_4\[23\] ci_neuron.uut_simple_neuron.titan_id_3\[23\]
+ _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04989_ _00689_ _00042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06728_ _01947_ _01988_ _02365_ _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09516_ _03851_ ci_neuron.input_memory\[1\]\[21\] _01368_ _02804_ _04716_ _04717_
+ _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_09447_ _04652_ _04670_ _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06659_ _02259_ _02298_ _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_66_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09378_ _04598_ _04601_ _04609_ _04612_ _00516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_47_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08329_ _03839_ _03842_ _03843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_35_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10222_ _00127_ net186 ci_neuron.uut_simple_neuron.titan_id_6\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10153_ _00218_ net236 ci_neuron.uut_simple_neuron.titan_id_3\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10084_ _00181_ net107 ci_neuron.uut_simple_neuron.titan_id_0\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07105__A2 _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07700_ ci_neuron.uut_simple_neuron.titan_id_4\[10\] ci_neuron.uut_simple_neuron.titan_id_3\[10\]
+ _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05961_ _01619_ _01531_ _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05892_ _01550_ _01552_ _01553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08680_ _04135_ _04141_ _04147_ _04148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_04912_ _00644_ _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07631_ _02132_ _03188_ _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04843_ internal_ih.current_instruction\[1\] _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07562_ _02542_ _02562_ _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06513_ _02077_ _02107_ _02156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09301_ _04545_ _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09341__I0 _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07493_ _02898_ _03050_ _03119_ _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_06444_ _01955_ _02052_ _02087_ _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09232_ _04499_ _04519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_118_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06375_ _02018_ _02019_ _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09163_ ci_neuron.uut_simple_neuron.titan_id_6\[25\] _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05326_ _00997_ _00998_ _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08114_ _03659_ _00073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09094_ _04415_ _04435_ _04436_ _00408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_102_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05257_ _00905_ _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_56_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08045_ ci_neuron.uut_simple_neuron.titan_id_1\[5\] ci_neuron.uut_simple_neuron.titan_id_0\[5\]
+ _03601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_116_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05188_ ci_neuron.uut_simple_neuron.x2\[6\] _00861_ _00866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09996_ _00511_ net92 ci_neuron.input_memory\[1\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08947_ internal_ih.byte6\[0\] internal_ih.byte5\[0\] _04317_ _04320_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08878_ internal_ih.byte2\[2\] internal_ih.byte1\[2\] _04280_ _04281_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07829_ ci_neuron.uut_simple_neuron.titan_id_2\[1\] ci_neuron.uut_simple_neuron.titan_id_5\[1\]
+ _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09332__I0 _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07271__A1 _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05821__A2 _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07023__A1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10205_ _00101_ net270 ci_neuron.uut_simple_neuron.titan_id_5\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08771__A1 _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10136_ _00201_ net274 ci_neuron.uut_simple_neuron.titan_id_3\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10142__D _00207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10067_ _00194_ net201 ci_neuron.uut_simple_neuron.titan_id_0\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08895__I _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09323__I0 _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06160_ _01767_ _01809_ _01814_ _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_124_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07262__A1 _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06091_ _01707_ _01708_ _01716_ _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05111_ _00791_ _00767_ _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05042_ _00727_ _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__08762__A1 _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09850_ _00429_ net158 ci_neuron.output_memory\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06993_ _02495_ _02626_ _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08801_ _04208_ _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09781_ _00360_ net47 internal_ih.byte3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05944_ _01255_ _01566_ _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08732_ _04185_ _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08663_ net5 _04131_ _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout67_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05875_ _01535_ _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07614_ ci_neuron.uut_simple_neuron.x3\[30\] _02611_ _03238_ _03239_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09314__I0 _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08594_ _04019_ _04071_ _04072_ _04073_ _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_48_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07545_ _02939_ _03170_ _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08817__A2 _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07476_ _02497_ _03102_ _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_64_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06427_ _02033_ _02063_ _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_62_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09215_ _04023_ _03795_ _04509_ _04510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06358_ _02000_ _02003_ _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_60_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09146_ _04469_ _00427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06289_ _01824_ _01936_ _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07253__A1 _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05309_ _00982_ _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06056__A2 _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09077_ _04405_ _04420_ _04421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08028_ ci_neuron.uut_simple_neuron.titan_id_1\[4\] ci_neuron.uut_simple_neuron.titan_id_0\[4\]
+ _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05567__A1 _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09979_ _00494_ net229 ci_neuron.input_memory\[1\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_129_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07547__A2 _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08595__I1 _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10119_ _00243_ net238 ci_neuron.uut_simple_neuron.titan_id_4\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout271_I net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05660_ _00859_ _01178_ _01324_ _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_77_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05591_ _01222_ _01229_ _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07330_ _02956_ _02958_ _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07261_ _02889_ _02818_ _02890_ _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07483__A1 _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09000_ _04349_ _00401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07192_ _01883_ _02755_ _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06212_ _01862_ _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06143_ _01749_ _01768_ _01797_ _01798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06074_ _01647_ _01685_ _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05025_ ci_neuron.instruction_i\[3\] ci_neuron.instruction_i\[5\] _00711_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09902_ _00021_ net14 ci_neuron.address_i\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09833_ _00412_ net158 ci_neuron.output_memory\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06976_ _02279_ _02561_ _02609_ _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09764_ _00343_ net60 internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05927_ _01527_ _01586_ _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08715_ internal_ih.spi_rx_byte_i\[3\] _04171_ _04175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09695_ net1 net57 spi_interface_cvonk.SCLK_r\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05858_ _01470_ _01485_ _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08646_ _04117_ _00279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_64_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05789_ _01450_ _01443_ _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05721__A1 _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08577_ _04059_ _02616_ _04053_ _04060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07528_ _03118_ _03132_ _03153_ _03154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07459_ _02934_ _03008_ _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09129_ ci_neuron.uut_simple_neuron.titan_id_6\[8\] _04461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_75_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08577__I1 _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06179__B _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout117_I net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07029__I _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06830_ _02256_ _02299_ _02354_ _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06761_ _02372_ _02398_ _02399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06692_ _02329_ _02330_ _02331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05712_ _01375_ _01337_ _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09480_ ci_neuron.output_memory\[16\] _04698_ _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08500_ _03945_ _03992_ _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05643_ _01247_ _01308_ _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08431_ _03929_ _03931_ _03932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05703__A1 _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05574_ _01166_ _01199_ _01201_ _01242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08362_ _03861_ ci_neuron.uut_simple_neuron.x0\[23\] _03871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07313_ _02932_ _02941_ _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08293_ _03796_ _03808_ _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07244_ _02548_ _02725_ _02874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07175_ _02804_ _02805_ _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06126_ _01779_ _01781_ _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06057_ _01710_ _01711_ _01713_ _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_2_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05008_ internal_ih.byte3\[3\] _00696_ _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_6_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09816_ _00395_ net58 internal_ih.current_instruction\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_126_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06959_ _01850_ _02592_ _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09747_ _00326_ net218 ci_neuron.uut_simple_neuron.x2\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09678_ _00265_ net232 ci_neuron.uut_simple_neuron.x3\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08629_ _03900_ _04102_ _04097_ _03892_ _03943_ _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__05170__A2 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07998__A2 ci_neuron.uut_simple_neuron.titan_id_5\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10150__D _00215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09427__A2 _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout234_I net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05290_ _00963_ _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_110_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08980_ internal_ih.byte7\[7\] internal_ih.byte6\[7\] _04257_ _04338_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07931_ _03506_ _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07862_ _03446_ _03447_ _03449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_3_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06813_ _02447_ _02449_ _02450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09601_ _04796_ _00555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07793_ _03390_ _03392_ _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09532_ _04696_ _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06744_ _02223_ _02340_ _02381_ _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_06675_ _02313_ _02274_ _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09463_ ci_neuron.output_val_internal\[13\] _04680_ _04685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_121_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05626_ _01289_ _01291_ _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04846__I _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09394_ ci_neuron.output_val_internal\[3\] _04611_ _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08414_ ci_neuron.uut_simple_neuron.x0\[30\] _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05557_ _01192_ _01224_ _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08345_ ci_neuron.uut_simple_neuron.x0\[21\] ci_neuron.uut_simple_neuron.x0\[22\]
+ _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_50_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05488_ _01124_ _01157_ _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08276_ ci_neuron.uut_simple_neuron.x0\[13\] _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07227_ _02811_ _02814_ _02856_ _02857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07158_ _02787_ _02788_ _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_100_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06109_ _01713_ _01763_ _01764_ _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07089_ _02678_ _02684_ _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_72_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout131 net132 net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout120 net121 net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout142 net145 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout164 net216 net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout153 net156 net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06301__I _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout175 net176 net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout197 net198 net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout186 net190 net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_69_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09432__I2 _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_94_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06159__A1 ci_neuron.uut_simple_neuron.x2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08943__I1 internal_ih.byte4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05906__A1 _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06460_ _02103_ _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_88_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05411_ _01048_ _01051_ _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06391_ _01987_ _02034_ _02035_ _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08130_ ci_neuron.uut_simple_neuron.titan_id_1\[21\] ci_neuron.uut_simple_neuron.titan_id_0\[21\]
+ _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05342_ _01013_ _01014_ _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06634__A2 _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05273_ _00946_ _00947_ _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08061_ _03607_ _03612_ _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07012_ _02641_ _02645_ _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout97_I net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08963_ internal_ih.byte6\[7\] internal_ih.byte5\[7\] _04327_ _04329_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07914_ _03489_ _03490_ _03492_ _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08894_ _04289_ _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07845_ ci_neuron.uut_simple_neuron.titan_id_2\[4\] ci_neuron.uut_simple_neuron.titan_id_5\[4\]
+ _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07776_ _03378_ _00110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06570__A1 _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04988_ internal_ih.byte2\[2\] _00686_ _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06727_ _01946_ _01952_ _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09515_ ci_neuron.output_memory\[21\] _04722_ _04729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09446_ _03783_ ci_neuron.input_memory\[1\]\[11\] _00977_ _02139_ _04667_ _04669_
+ _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_06658_ _02262_ _02297_ _02298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_82_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06589_ _02139_ _02187_ _02229_ _02230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05609_ _01251_ _01275_ _01276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09377_ ci_neuron.output_val_internal\[0\] _04611_ _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08328_ _03840_ _03841_ _03833_ _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07822__A1 ci_neuron.uut_simple_neuron.titan_id_4\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08259_ _03781_ _00170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06389__A1 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10221_ _00119_ net44 ci_neuron.uut_simple_neuron.titan_id_5\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10152_ _00217_ net237 ci_neuron.uut_simple_neuron.titan_id_3\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09327__A1 ci_neuron.input_memory\[1\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10083_ _00180_ net108 ci_neuron.uut_simple_neuron.titan_id_0\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_13_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08613__I0 _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05960_ ci_neuron.uut_simple_neuron.x2\[26\] _01619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05891_ _01493_ _01551_ _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04911_ internal_ih.byte5\[2\] _00640_ _00641_ internal_ih.byte1\[2\] _00644_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07630_ _02542_ _02562_ _03255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04842_ internal_ih.current_instruction\[0\] internal_ih.current_instruction\[1\]
+ internal_ih.current_instruction\[2\] _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_07561_ _03185_ _03186_ _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06512_ _02077_ _02107_ _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_105_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09300_ _04010_ _04546_ _04560_ _00490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07492_ _03047_ _03049_ _03119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_8_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06443_ _02085_ _02086_ _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_63_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09231_ _04518_ _00463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06374_ _02018_ _02019_ _02020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_17_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09162_ _04477_ _00435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05325_ _00962_ _00987_ _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08113_ _03657_ _03658_ _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_126_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08852__I0 internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09093_ internal_ih.spi_tx_byte_o\[5\] _04427_ _04436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05256_ _00907_ _00920_ _00931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08044_ _03600_ _00091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05187_ _00812_ _00846_ _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05291__A1 _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09995_ _00510_ net89 ci_neuron.input_memory\[1\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08946_ _04319_ _00377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08877_ _04269_ _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07828_ ci_neuron.uut_simple_neuron.titan_id_2\[0\] ci_neuron.uut_simple_neuron.titan_id_5\[0\]
+ _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07759_ ci_neuron.uut_simple_neuron.titan_id_4\[20\] ci_neuron.uut_simple_neuron.titan_id_3\[20\]
+ _03364_ _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_67_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09429_ ci_neuron.output_val_internal\[8\] _04655_ _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10204_ _00100_ net270 ci_neuron.uut_simple_neuron.titan_id_5\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10135_ _00227_ net273 ci_neuron.uut_simple_neuron.titan_id_3\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10066_ _00193_ net188 ci_neuron.uut_simple_neuron.titan_id_0\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout147_I net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05110_ _00773_ _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08834__I0 internal_ih.byte0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06090_ _01744_ _01745_ _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05041_ ci_neuron.address_i\[2\] _00726_ _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_0_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08800_ _04235_ _00315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06992_ _02622_ _02625_ _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09780_ _00359_ net50 internal_ih.byte3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05943_ _01557_ _01565_ _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08731_ _04173_ _04174_ _04181_ _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_56_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08662_ _04124_ _04126_ _04131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07613_ _01850_ _03228_ _03237_ _03238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_89_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05874_ _01528_ _01530_ _01534_ _01535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_88_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08593_ ci_neuron.value_i\[21\] _04013_ _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07544_ _03168_ _03169_ _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07475_ _02504_ _03101_ _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06426_ _02026_ _02068_ _02069_ _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_91_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09214_ _04499_ _04509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08326__I _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06357_ _01960_ _02002_ _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08825__I0 _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09145_ ci_neuron.uut_simple_neuron.titan_id_6\[16\] _04469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06288_ _01858_ _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05308_ _00981_ _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09076_ _04419_ ci_neuron.stream_o\[12\] _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05239_ _00912_ _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08027_ ci_neuron.uut_simple_neuron.titan_id_1\[4\] ci_neuron.uut_simple_neuron.titan_id_0\[4\]
+ _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09250__I0 _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09978_ _00493_ net229 ci_neuron.input_memory\[1\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08929_ _04309_ _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_129_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09241__I0 _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06755__A1 _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10118_ _00242_ net238 ci_neuron.uut_simple_neuron.titan_id_4\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10049_ _00534_ net138 ci_neuron.output_val_internal\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout264_I net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Left_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_102_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05590_ _01252_ _01219_ _01256_ _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07260_ _02326_ _02817_ _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07191_ _02217_ _02237_ _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06211_ _01823_ _01861_ _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08590__B _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06142_ _01700_ _01769_ _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06073_ _01682_ _01684_ _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_20_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09901_ _00020_ net11 ci_neuron.address_i\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05024_ _00708_ _00709_ _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_113_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09832_ _00411_ net153 ci_neuron.output_memory\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09763_ _00342_ net67 internal_ih.byte1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06975_ _02280_ _02441_ _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08714_ internal_ih.spi_rx_byte_i\[1\] internal_ih.spi_rx_byte_i\[0\] internal_ih.spi_rx_byte_i\[2\]
+ _04174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_05926_ _01576_ _01585_ _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09694_ _00281_ net92 ci_neuron.uut_simple_neuron.x3\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05857_ _01412_ _01516_ _01517_ _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08645_ _04116_ ci_neuron.uut_simple_neuron.x3\[29\] _04111_ _04117_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08576_ _04056_ _04058_ _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_124_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07527_ _03075_ _03117_ _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05788_ _01449_ _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07458_ _03083_ _03084_ _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06409_ _02047_ _02053_ _02054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07389_ _02676_ _02858_ _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09128_ _04460_ _00418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05237__A1 _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09059_ _04378_ _04403_ _04404_ _00405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08726__A2 _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06737__A1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07217__A2 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06728__A1 _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06760_ _02376_ _02378_ _02397_ _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06691_ _02286_ _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05711_ _01332_ _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05642_ _01076_ _01234_ _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_59_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08430_ ci_neuron.normalised_stream_write_address\[0\] _03930_ _03927_ _03931_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05573_ _01166_ _01199_ _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08361_ _03861_ _03863_ _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07312_ _02933_ _02940_ _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08292_ ci_neuron.uut_simple_neuron.x0\[15\] _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07243_ _02862_ _02872_ _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07174_ _02731_ _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06125_ _01731_ _01780_ _01728_ _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_41_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06056_ _01573_ _01579_ _01712_ _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05007_ _00699_ _00051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_6_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09815_ _00394_ net58 internal_ih.current_instruction\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_126_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06958_ _02590_ _02591_ _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09746_ _00325_ net218 ci_neuron.uut_simple_neuron.x2\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09677_ _00264_ net232 ci_neuron.uut_simple_neuron.x3\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05909_ _01530_ _01534_ _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06889_ _02524_ _00238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08628_ _03878_ _04081_ _04102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_77_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08559_ _04043_ _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08644__A1 _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05697__A1 _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07930_ ci_neuron.uut_simple_neuron.titan_id_2\[17\] ci_neuron.uut_simple_neuron.titan_id_5\[17\]
+ ci_neuron.uut_simple_neuron.titan_id_2\[16\] ci_neuron.uut_simple_neuron.titan_id_5\[16\]
+ _03506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_48_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07861_ _03448_ _00155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07792_ _03387_ _03388_ _03391_ _03392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06812_ _02383_ _02448_ _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09600_ ci_neuron.stream_o\[4\] ci_neuron.output_memory\[4\] _04795_ _04796_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06743_ _02379_ _02380_ _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_64_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09531_ _04721_ _04737_ _04741_ _04742_ _00539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__07126__A1 _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06674_ _01899_ _02313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_108_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09462_ _04677_ _04683_ _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05625_ _01227_ _01290_ _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09393_ _04603_ _04624_ _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08413_ _03905_ _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_121_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05556_ _01104_ _01223_ _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08535__S _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08344_ _03855_ _00181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_50_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05487_ _01126_ _01156_ _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06101__A2 _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08275_ _03794_ _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07226_ _02803_ _02810_ _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_89_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04862__I _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07157_ _01921_ _02313_ _02714_ _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__05860__A1 _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06108_ _01706_ _01667_ _01710_ _01764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07088_ _02688_ _02692_ _02719_ _02720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_72_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06039_ _01374_ _01659_ _01695_ _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout110 net111 net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout121 net122 net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07365__A1 _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout132 net134 net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout143 net145 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout154 net156 net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout165 net167 net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout176 net181 net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout198 net199 net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout187 net190 net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09729_ _00308_ net253 ci_neuron.uut_simple_neuron.x2\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05851__A1 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09432__I3 _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout177_I net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05410_ _01034_ _01079_ _01080_ _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_68_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06390_ _01993_ _02011_ _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05341_ _00980_ _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05272_ _00944_ _00945_ _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08060_ ci_neuron.uut_simple_neuron.titan_id_1\[9\] ci_neuron.uut_simple_neuron.titan_id_0\[9\]
+ _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07011_ _02642_ _02644_ _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08962_ _04328_ _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07913_ ci_neuron.uut_simple_neuron.titan_id_2\[14\] ci_neuron.uut_simple_neuron.titan_id_5\[14\]
+ _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08893_ internal_ih.byte3\[1\] internal_ih.byte2\[1\] _04285_ _04289_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07844_ _03431_ _03433_ _03434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_3_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07775_ _03376_ _03377_ _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04987_ _00688_ _00041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06726_ _02362_ _02363_ _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_69_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04857__I _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09514_ _04721_ _04723_ _04726_ _04728_ _00536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06657_ _02268_ _02296_ _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07233__I ci_neuron.uut_simple_neuron.x3\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09445_ _04668_ _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05608_ _01257_ _01274_ _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06588_ _02226_ _02228_ _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09376_ _04610_ _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05539_ _01177_ _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08327_ _03835_ _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08258_ _03777_ _03780_ _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_50_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_49_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07209_ _02779_ _02839_ _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08189_ ci_neuron.uut_simple_neuron.titan_id_1\[31\] ci_neuron.uut_simple_neuron.titan_id_0\[31\]
+ _03721_ _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_10220_ _00117_ net45 ci_neuron.uut_simple_neuron.titan_id_5\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10151_ _00216_ net237 ci_neuron.uut_simple_neuron.titan_id_3\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05061__A2 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10082_ _00179_ net114 ci_neuron.uut_simple_neuron.titan_id_0\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_58_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_67_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08613__I1 _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07329__A1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04910_ _00643_ _00024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09680__D _00267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05890_ _01500_ _01502_ _01508_ _01495_ _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_45_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04841_ internal_ih.current_instruction\[5\] internal_ih.current_instruction\[4\]
+ internal_ih.current_instruction\[7\] internal_ih.current_instruction\[6\] _00592_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_07560_ _02497_ _03102_ _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06511_ _02122_ _02153_ _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_105_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07491_ _03075_ _03117_ _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09230_ _04064_ _03852_ _04514_ _04518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06442_ _02051_ _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06373_ _01975_ _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09161_ ci_neuron.uut_simple_neuron.titan_id_6\[24\] _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05324_ _00966_ _00986_ _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08112_ ci_neuron.uut_simple_neuron.titan_id_1\[18\] ci_neuron.uut_simple_neuron.titan_id_0\[18\]
+ _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09092_ ci_neuron.stream_o\[29\] _04416_ _04434_ _04435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08043_ _03598_ _03599_ _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05255_ _00930_ _00201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05186_ _00863_ _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09994_ _00509_ net89 ci_neuron.input_memory\[1\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08945_ internal_ih.byte5\[7\] internal_ih.byte4\[7\] _04317_ _04319_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09443__I _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08876_ _04279_ _00347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07827_ _03420_ _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07758_ _03360_ _03362_ _03363_ _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06709_ _02321_ _02347_ _02348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_80_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07689_ _03306_ _00124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09428_ _04610_ _04655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09359_ _04373_ _04593_ _04594_ _00515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_124_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05806__A1 _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08843__I1 _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07559__A1 _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09548__A2 _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10203_ _00099_ net278 ci_neuron.uut_simple_neuron.titan_id_5\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10134_ _00226_ net273 ci_neuron.uut_simple_neuron.titan_id_3\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10065_ _00190_ net187 ci_neuron.uut_simple_neuron.titan_id_0\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_75_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08834__I1 _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05040_ _00722_ _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_84_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09003__A4 _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06991_ _02551_ _02624_ _02625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05942_ _01560_ _01590_ _01600_ _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08730_ internal_ih.received_byte_count\[1\] _04189_ _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05873_ _00739_ _01531_ _01533_ _01474_ _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_08661_ _04124_ _04126_ _04129_ _04130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07612_ _02802_ _03233_ _03236_ _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_89_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08592_ _03848_ _03850_ _04066_ _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_07543_ ci_neuron.uut_simple_neuron.x3\[29\] _03088_ _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_93_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07474_ _02812_ _03019_ _03018_ _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06425_ _02066_ _02067_ _02064_ _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_57_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09213_ _03785_ _04489_ _04508_ _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09144_ _04468_ _00426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06356_ ci_neuron.uut_simple_neuron.x3\[8\] _02001_ _02002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06287_ _01860_ _01934_ _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_05307_ _00866_ _00976_ _00980_ _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09075_ _04361_ _04419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05238_ _00895_ _00911_ _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08026_ _03585_ _00088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05169_ _00846_ _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_12_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08202__A2 _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09977_ _00492_ net174 ci_neuron.input_memory\[1\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08928_ internal_ih.byte5\[0\] internal_ih.byte4\[0\] _04306_ _04309_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_129_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08859_ _04269_ _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_79_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09927__CLK net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10117_ _00241_ net245 ci_neuron.uut_simple_neuron.titan_id_4\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10048_ _00533_ net138 ci_neuron.output_val_internal\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06210_ _01858_ _01860_ _01861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07190_ _02794_ _02820_ _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_115_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06141_ _01754_ _01794_ _01795_ _01796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06072_ _01727_ _01728_ _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09900_ _00019_ net11 ci_neuron.address_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05023_ ci_neuron.instruction_i\[1\] _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09831_ _00410_ net126 internal_ih.spi_tx_byte_o\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06974_ _02544_ _02565_ _02607_ _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08991__I0 _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09762_ _00341_ net60 internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout72_I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06410__I _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05925_ _01530_ _01584_ _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08713_ _04170_ internal_ih.spi_rx_byte_i\[3\] _04172_ _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_83_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09693_ _00280_ net90 ci_neuron.uut_simple_neuron.x3\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05856_ _01413_ _01466_ _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08644_ _04019_ _04113_ _04114_ _04115_ _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_95_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05787_ _01124_ _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08575_ _03841_ _04044_ _04057_ _03943_ _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_124_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07526_ _03120_ _03131_ _03151_ _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07457_ ci_neuron.uut_simple_neuron.x3\[27\] _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07388_ _03011_ _03015_ _03016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06408_ _01955_ _02052_ _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06339_ _01847_ _01984_ _01985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_20_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08423__A2 _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09127_ ci_neuron.uut_simple_neuron.titan_id_6\[7\] _04460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05237__A2 _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09058_ internal_ih.spi_tx_byte_o\[2\] _04379_ _04404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08009_ _03569_ _03571_ _03572_ _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06737__A2 _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06673__A1 _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06690_ _02285_ _02329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05710_ _01371_ _01373_ _01374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05641_ _01243_ _01305_ _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08360_ ci_neuron.uut_simple_neuron.x0\[23\] ci_neuron.uut_simple_neuron.x0\[24\]
+ _03869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07311_ _02936_ _02939_ _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05572_ _01235_ _01239_ _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__04911__B2 internal_ih.byte1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08291_ _03808_ _03809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07242_ _02682_ _02871_ _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_27_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07173_ _02734_ _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06124_ _01682_ _01684_ _01727_ _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06055_ _01473_ _01577_ _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10074__D _00171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04978__A1 internal_ih.byte1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05006_ internal_ih.byte3\[2\] _00696_ _00699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09814_ _00393_ net40 internal_ih.byte7\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_126_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06957_ _02531_ _02537_ _02591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09745_ _00324_ net218 ci_neuron.uut_simple_neuron.x2\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06888_ _02521_ _02523_ _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09676_ _00263_ net232 ci_neuron.uut_simple_neuron.x3\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05908_ _01567_ _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05839_ _01498_ _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08627_ ci_neuron.value_i\[27\] _04055_ _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_25_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08558_ _03821_ _04038_ _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__04902__B2 internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04902__A1 internal_ih.byte4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07509_ _02996_ _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_65_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08489_ ci_neuron.value_i\[6\] _03944_ _03983_ _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_91_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__04969__A1 internal_ih.byte1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09626__I _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07860_ _03446_ _03447_ _03448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07791_ ci_neuron.uut_simple_neuron.titan_id_4\[25\] ci_neuron.uut_simple_neuron.titan_id_3\[25\]
+ _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06811_ ci_neuron.uut_simple_neuron.x3\[17\] ci_neuron.uut_simple_neuron.x3\[18\]
+ _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_3_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06742_ _02339_ _02380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09530_ ci_neuron.output_val_internal\[23\] _04727_ _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09461_ _03797_ ci_neuron.input_memory\[1\]\[13\] _01006_ _02228_ _04667_ _04669_
+ _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_06673_ _01908_ _02273_ _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05624_ ci_neuron.uut_simple_neuron.x2\[19\] ci_neuron.uut_simple_neuron.x2\[20\]
+ _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09392_ _03730_ ci_neuron.input_memory\[1\]\[3\] _00758_ _01872_ _04622_ _04623_
+ _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_59_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout35_I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08412_ _03914_ _00191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_121_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05555_ _01096_ _01149_ _01184_ _01223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08343_ _03849_ _03851_ _03854_ _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_50_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08274_ ci_neuron.uut_simple_neuron.x0\[12\] _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07225_ _02796_ _02853_ _02854_ _02815_ _02819_ _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_05486_ _01130_ _01134_ _01155_ _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_73_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07156_ _02785_ _02786_ _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07087_ _02675_ _02687_ _02719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06107_ _01578_ _01711_ _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_30_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06038_ _01462_ _01660_ _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_72_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout111 net116 net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout122 net127 net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout100 net101 net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout133 net134 net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout144 net145 net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout155 net157 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05376__A1 _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout177 net180 net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout166 net167 net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout199 net214 net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout188 net189 net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09728_ _00307_ net254 ci_neuron.uut_simple_neuron.x2\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07989_ _03551_ _03552_ _03555_ _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09181__I _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09659_ ci_neuron.stream_o\[30\] ci_neuron.output_memory\[30\] _04826_ _04829_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09290__A2 _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06800__A1 _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08928__I0 internal_ih.byte5\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07604__I _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05340_ _00811_ _00861_ _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09281__A2 _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05271_ _00944_ _00945_ _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07010_ _02573_ _02643_ _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08961_ internal_ih.byte6\[6\] internal_ih.byte5\[6\] _04327_ _04328_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07912_ _03491_ _00132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08892_ _04288_ _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07843_ _03429_ _03432_ _03433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07774_ ci_neuron.uut_simple_neuron.titan_id_4\[23\] ci_neuron.uut_simple_neuron.titan_id_3\[23\]
+ _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04986_ internal_ih.byte2\[1\] _00686_ _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06725_ _01929_ _02324_ _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09513_ ci_neuron.output_val_internal\[20\] _04727_ _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06656_ _02271_ _02295_ _02296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09444_ _03935_ _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05607_ _01259_ _01273_ _01274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06587_ _02227_ _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05530__A1 _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09375_ _04596_ _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05538_ _01170_ _01196_ _01205_ _01206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08326_ _03824_ _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05469_ _01042_ _01093_ _01138_ _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08257_ _03778_ _03779_ _03780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07208_ _02835_ _02838_ _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_104_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_104_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08188_ _03717_ _03718_ _03720_ _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07139_ _02770_ _00242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07035__A1 _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09176__I _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10150_ _00215_ net239 ci_neuron.uut_simple_neuron.titan_id_3\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10081_ _00178_ net114 ci_neuron.uut_simple_neuron.titan_id_0\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09583__I0 _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_113_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_122_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_13_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08774__A1 _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10279_ _00572_ net183 ci_neuron.stream_o\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_04840_ _00591_ internal_ih.got_all_data vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07490_ _03106_ _03116_ _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06510_ _02124_ _02152_ _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_105_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06441_ _02049_ _02085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06372_ _01972_ _02018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09160_ _04476_ _00434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05323_ _00959_ _00989_ _00995_ _00996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08111_ _03652_ _03654_ _03656_ _03657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09091_ _04356_ _04431_ _04433_ _04411_ _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_44_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05254_ _00926_ _00929_ _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08042_ ci_neuron.uut_simple_neuron.titan_id_1\[7\] ci_neuron.uut_simple_neuron.titan_id_0\[7\]
+ _03599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05185_ _00781_ _00838_ _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08765__A1 _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09993_ _00508_ net89 ci_neuron.input_memory\[1\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08944_ _04318_ _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08875_ internal_ih.byte2\[1\] internal_ih.byte1\[1\] _04275_ _04279_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07826_ ci_neuron.uut_simple_neuron.titan_id_4\[1\] ci_neuron.uut_simple_neuron.titan_id_3\[1\]
+ _03420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07757_ ci_neuron.uut_simple_neuron.titan_id_4\[19\] ci_neuron.uut_simple_neuron.titan_id_3\[19\]
+ _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_04969_ internal_ih.byte1\[2\] _00675_ _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06708_ _02325_ _02328_ _02346_ _02347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_67_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07688_ _03304_ _03305_ _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06639_ _02230_ _02279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_80_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09427_ _04652_ _04653_ _04654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_81_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09358_ _04385_ _04373_ _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07256__A1 _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08309_ _03810_ _03825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_10_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09289_ _03979_ _04553_ _04554_ _00485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10202_ _00098_ net278 ci_neuron.uut_simple_neuron.titan_id_5\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10133_ _00225_ net273 ci_neuron.uut_simple_neuron.titan_id_3\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10064_ _00065_ net189 ci_neuron.uut_simple_neuron.titan_id_0\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09308__I0 _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09484__A2 _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07495__A1 _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06298__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05402__I _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06990_ ci_neuron.uut_simple_neuron.x3\[20\] _02623_ _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05941_ _01563_ _01589_ _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05872_ _01475_ _01532_ _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08660_ spi_interface_cvonk.buffer\[7\] internal_ih.spi_tx_byte_o\[7\] _04128_ _04129_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07611_ _03234_ _03235_ _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08591_ _03849_ _04066_ _03851_ _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07542_ _03166_ _03167_ _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07486__A1 _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07473_ _03099_ _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06424_ _02066_ _02067_ _02064_ _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09212_ _04017_ _04496_ _04508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06355_ ci_neuron.uut_simple_neuron.x3\[9\] _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09143_ ci_neuron.uut_simple_neuron.titan_id_6\[15\] _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_118_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05306_ _00895_ _00978_ _00979_ _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06286_ _01931_ _01933_ _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09074_ _04359_ _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_97_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05237_ _00750_ _00896_ _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08025_ ci_neuron.uut_simple_neuron.titan_id_1\[4\] ci_neuron.uut_simple_neuron.titan_id_0\[4\]
+ _03584_ _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_4_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05168_ ci_neuron.uut_simple_neuron.x2\[7\] _00846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07410__A1 _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05099_ _00742_ _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09976_ _00491_ net253 ci_neuron.input_memory\[1\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09454__I _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08927_ _04308_ _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_129_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08858_ _04256_ _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_129_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07809_ _03391_ _03394_ _03405_ _03406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08789_ _04229_ _00310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05378__B _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10236__CLK net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07401__A1 _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10116_ _00240_ net245 ci_neuron.uut_simple_neuron.titan_id_4\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10047_ _00532_ net166 ci_neuron.output_val_internal\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout152_I net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06140_ _01792_ _01793_ _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08443__I _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06071_ _01687_ _01688_ _01726_ _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_111_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05022_ ci_neuron.instruction_i\[0\] _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_113_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08599__B _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09274__I _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09830_ _00409_ net139 internal_ih.spi_tx_byte_o\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06973_ _02546_ _02564_ _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05508__S _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09761_ _00340_ net70 internal_ih.byte1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05924_ _01577_ _01581_ _01583_ _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08712_ internal_ih.spi_rx_byte_i\[1\] _04143_ _04171_ _04172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09692_ _00279_ net90 ci_neuron.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_05855_ _01413_ _01466_ _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08643_ ci_neuron.value_i\[29\] _04013_ _04115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05786_ _01411_ _01442_ _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08574_ _03832_ _04043_ _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_124_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07525_ _03123_ _03130_ _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07459__A1 _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07456_ _02937_ _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_92_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06682__A2 _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07387_ _03013_ _02939_ _03014_ _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06407_ _02049_ _02051_ _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_79_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06338_ _01983_ _01984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09126_ _04459_ _00417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06269_ _01909_ _01911_ _01917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09057_ ci_neuron.stream_o\[26\] _04381_ _04402_ _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08008_ ci_neuron.uut_simple_neuron.titan_id_2\[29\] ci_neuron.uut_simple_neuron.titan_id_5\[29\]
+ _03572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06198__A1 _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09384__A1 ci_neuron.output_memory\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09959_ _00474_ net74 ci_neuron.uut_simple_neuron.x0\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09184__I _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05173__A2 _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06673__A2 _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07622__A1 _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05640_ _01244_ _01305_ _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08438__I _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05571_ _01236_ _01237_ _01238_ _01239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_63_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07310_ _02863_ _02938_ _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_86_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08290_ ci_neuron.uut_simple_neuron.x0\[14\] _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07241_ _02867_ _02870_ _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07172_ _02676_ _02802_ _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07613__A1 _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06123_ _01737_ _01778_ _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06054_ _01706_ _01667_ _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05005_ _00698_ _00050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09813_ _00392_ net40 internal_ih.byte7\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06956_ _02534_ _02536_ _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09744_ _00323_ net91 ci_neuron.uut_simple_neuron.x2\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_126_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06887_ _02466_ _02468_ _02522_ _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09675_ _00262_ net261 ci_neuron.uut_simple_neuron.x3\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05907_ _01254_ _01566_ _01567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05838_ _01123_ _01499_ _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08626_ _04100_ _00276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05769_ _01428_ _01429_ _01431_ _01432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_76_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_53_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08557_ _03822_ _04038_ _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07508_ _03071_ _03134_ _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08488_ _03945_ _03982_ _03983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07439_ _02778_ _02980_ _03062_ _03065_ _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__06655__A2 _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09109_ _04356_ _04447_ _04449_ _04370_ _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_103_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08891__I0 internal_ih.byte3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout115_I net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07790_ ci_neuron.uut_simple_neuron.titan_id_4\[26\] ci_neuron.uut_simple_neuron.titan_id_3\[26\]
+ _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06810_ _02333_ _02389_ _02446_ _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06741_ _02337_ _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09552__I _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09520__A1 ci_neuron.output_memory\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09460_ ci_neuron.output_memory\[13\] _04675_ _04682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06672_ _02268_ _02296_ _02310_ _02311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_108_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08411_ _03910_ _03913_ _03914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05623_ _00747_ _01268_ _01289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09391_ _04606_ _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_129_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05554_ _00742_ _01193_ _01222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08342_ _03852_ _03849_ _03853_ _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_50_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04896__B2 internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05485_ _01144_ _01154_ _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08273_ _03793_ _00172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07224_ _02811_ _02814_ _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07155_ _02751_ _02757_ _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07086_ _02668_ _02694_ _02717_ _02718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06106_ _01753_ _01761_ _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06037_ _01692_ _01693_ _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout112 net115 net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout101 net106 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout123 net125 net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout134 net135 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout145 net146 net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout156 net157 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout178 net180 net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07988_ ci_neuron.uut_simple_neuron.titan_id_2\[26\] ci_neuron.uut_simple_neuron.titan_id_5\[26\]
+ _03555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout167 net168 net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout189 net190 net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06939_ _02515_ _02517_ _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09727_ _00306_ net255 ci_neuron.uut_simple_neuron.x2\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06325__A1 _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09658_ _04828_ _00580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08609_ _04085_ _02928_ _04086_ _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09589_ _03926_ _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08873__I0 internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08625__I0 _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06800__A2 _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08928__I1 internal_ih.byte4\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08553__A2 _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09372__I _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06316__A1 _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout232_I net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08864__I0 internal_ih.byte1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05270_ _00751_ _00942_ _00918_ _00909_ _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_71_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08652__S _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08960_ _04311_ _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07911_ _03489_ _03490_ _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08919__I1 internal_ih.byte3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08891_ internal_ih.byte3\[0\] internal_ih.byte2\[0\] _04285_ _04288_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07842_ ci_neuron.uut_simple_neuron.titan_id_2\[3\] ci_neuron.uut_simple_neuron.titan_id_5\[3\]
+ _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07773_ _03372_ _03374_ _03375_ _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09512_ _04704_ _04727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04985_ _00687_ _00040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06724_ _01948_ _02323_ _02362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06655_ _02275_ _02294_ _02295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09443_ _04666_ _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_35_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05606_ _01261_ _01272_ _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09374_ _04603_ _04608_ _04609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06586_ ci_neuron.uut_simple_neuron.x3\[13\] _02227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08325_ _03837_ _03838_ _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05537_ _01172_ _01195_ _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_35_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05468_ _00983_ _01092_ _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08256_ _03755_ _03771_ ci_neuron.uut_simple_neuron.x0\[8\] _03779_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_6_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07207_ _02707_ _02836_ _02837_ _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08187_ ci_neuron.uut_simple_neuron.titan_id_1\[30\] ci_neuron.uut_simple_neuron.titan_id_0\[30\]
+ _03720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07138_ _02764_ _02766_ _02769_ _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_05399_ _01029_ _01027_ _01070_ _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07069_ _02638_ _02573_ _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_112_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10080_ _00177_ net113 ci_neuron.uut_simple_neuron.titan_id_0\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09192__I _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06849__A2 _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08472__S _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10278_ _00571_ net184 ci_neuron.stream_o\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08526__A2 _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06537__A1 _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout182_I net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06440_ _02054_ _02058_ _02083_ _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_105_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06371_ _01945_ _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05322_ _00946_ _00988_ _00995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08110_ ci_neuron.uut_simple_neuron.titan_id_1\[17\] ci_neuron.uut_simple_neuron.titan_id_0\[17\]
+ _03656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09090_ _04365_ _04432_ _04433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08462__A1 ci_neuron.value_i\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05253_ _00927_ _00928_ _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08041_ _03596_ _03597_ _03598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05184_ _00857_ _00860_ _00861_ _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_24_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09992_ _00507_ net85 ci_neuron.input_memory\[1\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout95_I net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08943_ internal_ih.byte5\[6\] internal_ih.byte4\[6\] _04317_ _04318_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08874_ _04278_ _00346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07825_ _03419_ _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07756_ ci_neuron.uut_simple_neuron.titan_id_4\[19\] ci_neuron.uut_simple_neuron.titan_id_3\[19\]
+ _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_04968_ _00677_ _00064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06707_ _02342_ _02345_ _02346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07687_ ci_neuron.uut_simple_neuron.titan_id_4\[8\] ci_neuron.uut_simple_neuron.titan_id_3\[8\]
+ _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09426_ _03770_ ci_neuron.input_memory\[1\]\[8\] _00867_ _01998_ _04644_ _04645_
+ _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_04899_ _00636_ _00020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09493__A3 _04709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06638_ _02235_ _02238_ _02277_ _02278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06569_ _01863_ _02175_ _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09357_ _04354_ _04592_ _04376_ _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09288_ ci_neuron.input_memory\[1\]\[5\] _04549_ _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08308_ _03823_ _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_10_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08239_ _03762_ _03763_ _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_35_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10201_ _00097_ net270 ci_neuron.uut_simple_neuron.titan_id_5\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10132_ _00224_ net266 ci_neuron.uut_simple_neuron.titan_id_3\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10063_ ci_neuron.uut_simple_neuron.x0\[0\] net183 ci_neuron.uut_simple_neuron.titan_id_0\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07192__A1 _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08819__I0 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05258__A1 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09244__I0 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05940_ _01599_ _00217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09547__I1 ci_neuron.input_memory\[1\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05871_ ci_neuron.uut_simple_neuron.x2\[25\] _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07610_ _02939_ _03170_ _03235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08590_ _02726_ _03941_ _04070_ _00270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07541_ _03084_ ci_neuron.uut_simple_neuron.x3\[28\] _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07472_ _03080_ _03098_ _03099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06423_ _02016_ _02022_ _02067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09211_ _04010_ _04503_ _04507_ _00454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06354_ _01959_ _01965_ _01999_ _02000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09142_ _04467_ _00425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05305_ _00910_ _00977_ _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_114_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06285_ _01878_ _01932_ _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09073_ _04361_ _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05236_ _00895_ _00911_ _00912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09235__I0 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08024_ _03580_ _03582_ _03583_ _03584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_102_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05167_ _00845_ _00225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_77_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05098_ _00763_ _00771_ _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09975_ _00490_ net175 ci_neuron.input_memory\[1\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08926_ internal_ih.byte4\[7\] internal_ih.byte3\[7\] _04306_ _04308_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_129_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08857_ _04268_ _00339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_129_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07808_ ci_neuron.uut_simple_neuron.titan_id_4\[26\] ci_neuron.uut_simple_neuron.titan_id_3\[26\]
+ _03405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06921__A1 ci_neuron.uut_simple_neuron.x3\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08788_ _04023_ _00971_ _04225_ _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07739_ ci_neuron.uut_simple_neuron.titan_id_4\[17\] ci_neuron.uut_simple_neuron.titan_id_3\[17\]
+ _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05488__A1 _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09409_ _04627_ _04635_ _04637_ _04638_ _00521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_125_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06988__A1 _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09226__I0 _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10115_ _00239_ net245 ci_neuron.uut_simple_neuron.titan_id_4\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10046_ _00531_ net166 ci_neuron.output_val_internal\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06979__A1 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06070_ _01687_ _01688_ _01726_ _01727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09217__I0 _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05021_ _00707_ _00065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_113_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09393__A2 _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06972_ _02599_ _02605_ _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09760_ _00339_ net67 internal_ih.byte1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05923_ _00738_ _01582_ _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09691_ _00278_ net218 ci_neuron.uut_simple_neuron.x3\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08711_ internal_ih.spi_rx_byte_i\[7\] internal_ih.spi_rx_byte_i\[6\] internal_ih.spi_rx_byte_i\[5\]
+ internal_ih.spi_rx_byte_i\[4\] _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_83_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08642_ _03900_ _03912_ _04102_ _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_05854_ _01513_ _01514_ _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05785_ _01447_ _00214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08573_ ci_neuron.value_i\[18\] _04055_ _04056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_124_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07524_ _03148_ _03149_ _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07455_ _02859_ _03010_ _03081_ _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06406_ _01964_ _02050_ _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_9_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07386_ _02933_ _02940_ _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06337_ _01830_ _01877_ _01982_ _01983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05890__A1 _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09125_ ci_neuron.uut_simple_neuron.titan_id_6\[6\] _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06268_ _01912_ _01914_ _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09056_ _04382_ _04399_ _04401_ _04354_ _04402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09208__I0 _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05642__A1 _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05219_ _00895_ _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08007_ ci_neuron.uut_simple_neuron.titan_id_2\[29\] ci_neuron.uut_simple_neuron.titan_id_5\[29\]
+ _03571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06199_ _01836_ _01839_ _01846_ _01850_ _00164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06198__A2 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09958_ _00473_ net76 ci_neuron.uut_simple_neuron.x0\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08909_ _04298_ _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07147__A1 _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09889_ _00050_ net21 ci_neuron.value_i\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_28_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05881__A1 _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_128_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09375__I _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10029_ ci_neuron.input_memory\[1\]\[29\] net86 ci_neuron.uut_simple_neuron.titan_id_1\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout262_I net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05570_ _01169_ _01197_ _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_63_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07240_ _02797_ _02869_ _02870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_73_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__04982__I _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07171_ _02799_ _02801_ _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05872__A1 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06122_ _01594_ _01777_ _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06053_ _01473_ _01577_ _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05004_ internal_ih.byte3\[1\] _00696_ _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09812_ _00391_ net39 internal_ih.byte7\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06955_ _02589_ _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09743_ _00322_ net219 ci_neuron.uut_simple_neuron.x2\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_126_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06886_ _02408_ _02406_ _02463_ _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09674_ _00261_ net261 ci_neuron.uut_simple_neuron.x3\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05906_ _01179_ _01565_ _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05837_ _01496_ _01305_ _01498_ _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08625_ _04099_ _03083_ _04086_ _04100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08556_ _04041_ _00265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07507_ _03073_ _03133_ _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05768_ _01344_ _01430_ _01431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_76_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05699_ _01341_ _01346_ _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_53_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08487_ _03753_ _03976_ _03982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07438_ _03059_ _03063_ _03064_ _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07369_ _02924_ _02949_ _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09108_ _04365_ _04448_ _04449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09039_ _04358_ ci_neuron.stream_o\[9\] _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06040__A1 _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09380__I2 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07540__A1 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08891__I1 internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10191__D _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06740_ _02342_ _02345_ _02377_ _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06671_ _02271_ _02295_ _02310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_108_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05622_ _00750_ _01287_ _01270_ _01263_ _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_08410_ _03907_ _03911_ _03912_ _03906_ _03913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_93_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09390_ _04604_ _04622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_121_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05553_ _01218_ _01220_ _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08341_ _03844_ _03846_ _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05484_ _01153_ _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08272_ _03789_ _03792_ _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_50_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07223_ _02811_ _02814_ _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_55_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08882__I1 internal_ih.byte1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09426__I3 _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07598__A1 _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07154_ _02754_ _02756_ _02785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09587__A2 _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07085_ _02671_ _02693_ _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06105_ _01714_ _01760_ _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06270__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06036_ _01568_ _01677_ _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout113 net115 net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout102 net104 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05048__I net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout124 net125 net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout135 net147 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout146 net147 net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout179 net180 net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout157 net162 net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07987_ ci_neuron.uut_simple_neuron.titan_id_2\[27\] ci_neuron.uut_simple_neuron.titan_id_5\[27\]
+ _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xfanout168 net172 net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06938_ _02569_ _02572_ _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_87_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09726_ _00305_ net255 ci_neuron.uut_simple_neuron.x2\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_2_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09511__A2 _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06869_ _02497_ _02504_ _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08570__I0 _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09657_ ci_neuron.stream_o\[29\] ci_neuron.output_memory\[29\] _04826_ _04828_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08608_ _03939_ _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09588_ _00710_ _00713_ _00725_ _04788_ _00550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_65_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08539_ ci_neuron.value_i\[13\] _04025_ _04026_ _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08873__I1 internal_ih.byte1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_98_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08625__I1 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06013__A1 _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08002__A2 ci_neuron.uut_simple_neuron.titan_id_5\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08864__I1 internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout225_I net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08732__I _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09569__A2 _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07910_ ci_neuron.uut_simple_neuron.titan_id_2\[14\] ci_neuron.uut_simple_neuron.titan_id_5\[14\]
+ _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08890_ _04287_ _00353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07841_ ci_neuron.uut_simple_neuron.titan_id_2\[3\] ci_neuron.uut_simple_neuron.titan_id_5\[3\]
+ _03431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07772_ ci_neuron.uut_simple_neuron.titan_id_4\[22\] ci_neuron.uut_simple_neuron.titan_id_3\[22\]
+ _03375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06723_ _02319_ _02348_ _02360_ _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_79_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04984_ internal_ih.byte2\[0\] _00686_ _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09511_ _04724_ _04725_ _04726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_69_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06654_ _02278_ _02293_ _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_91_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ _03930_ _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_35_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06585_ _02142_ _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_82_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05605_ _01262_ _01271_ _01272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09373_ _03725_ ci_neuron.input_memory\[1\]\[0\] _00736_ _02898_ _04605_ _04607_
+ _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_19_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05536_ _01204_ _00208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08324_ _03835_ ci_neuron.uut_simple_neuron.x0\[19\] _03838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10096__D _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05467_ _01083_ _01135_ _01136_ _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08255_ ci_neuron.uut_simple_neuron.x0\[8\] ci_neuron.uut_simple_neuron.x0\[9\] _03761_
+ _03764_ _03765_ _03778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_34_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07206_ _02709_ _02760_ _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05398_ _01065_ _01069_ _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08186_ _03719_ _00086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07137_ _02767_ _02768_ _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_18_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07068_ _02576_ _02641_ _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_93_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06019_ _01657_ _01676_ _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09709_ _00288_ net123 internal_ih.spi_rx_byte_i\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_27_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05809__A1 _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10277_ _00570_ net142 ci_neuron.stream_o\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06537__A2 _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08782__I0 _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_105_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06370_ _02015_ _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05321_ _00953_ _00956_ _00991_ _00951_ _00994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05252_ _00851_ _00875_ _00882_ _00902_ _00877_ _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_08040_ _03593_ _03594_ _03597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_54_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06225__A1 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05183_ ci_neuron.uut_simple_neuron.x2\[7\] ci_neuron.uut_simple_neuron.x2\[8\] _00861_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_116_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09991_ _00506_ net87 ci_neuron.input_memory\[1\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08942_ _04311_ _04317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_86_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08873_ internal_ih.byte2\[0\] internal_ih.byte1\[0\] _04275_ _04278_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07824_ ci_neuron.uut_simple_neuron.titan_id_4\[31\] ci_neuron.uut_simple_neuron.titan_id_3\[31\]
+ _03418_ _03419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_79_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07755_ _03361_ _00105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04967_ internal_ih.byte1\[1\] _00675_ _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06706_ _02344_ _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07686_ _03302_ _03303_ _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06637_ _02225_ _02276_ _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04898_ internal_ih.byte4\[5\] _00633_ _00634_ internal_ih.byte0\[5\] _00636_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09425_ _04602_ _04652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06568_ _02203_ _02205_ _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_81_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09356_ _04145_ _04179_ _04385_ _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06499_ ci_neuron.uut_simple_neuron.x3\[12\] _02142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05519_ _01186_ _01187_ _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_09287_ _04543_ _04553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08307_ ci_neuron.uut_simple_neuron.x0\[17\] _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_10_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08238_ _03752_ ci_neuron.uut_simple_neuron.x0\[7\] _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10200_ _00126_ net277 ci_neuron.uut_simple_neuron.titan_id_5\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08169_ ci_neuron.uut_simple_neuron.titan_id_1\[28\] ci_neuron.uut_simple_neuron.titan_id_0\[28\]
+ _03705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10131_ _00223_ net266 ci_neuron.uut_simple_neuron.titan_id_3\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10062_ _00547_ net167 ci_neuron.output_val_internal\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08819__I1 _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09547__I2 _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05870_ ci_neuron.uut_simple_neuron.x2\[24\] ci_neuron.uut_simple_neuron.x2\[25\]
+ _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07540_ _03083_ _03088_ _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07471_ _03093_ _03097_ _03098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06422_ _01981_ _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09210_ _04005_ _04496_ _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06353_ _01960_ _01998_ _01999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_84_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09141_ ci_neuron.uut_simple_neuron.titan_id_6\[14\] _04467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05304_ _00910_ _00977_ _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09072_ _04370_ _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06284_ ci_neuron.uut_simple_neuron.x3\[6\] ci_neuron.uut_simple_neuron.x3\[7\] _01932_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08023_ ci_neuron.uut_simple_neuron.titan_id_1\[3\] ci_neuron.uut_simple_neuron.titan_id_0\[3\]
+ _03583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05235_ _00910_ _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05166_ _00830_ _00831_ _00844_ _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_77_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05097_ _00736_ _00774_ _00772_ _00775_ _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XPHY_EDGE_ROW_71_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09974_ _00489_ net175 ci_neuron.input_memory\[1\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08925_ _04307_ _00368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05056__I _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08856_ internal_ih.byte1\[1\] internal_ih.byte0\[1\] _04264_ _04268_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_129_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07807_ _03390_ _03403_ _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05999_ _01655_ _01656_ _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08787_ _04228_ _00309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07738_ _03345_ _03346_ _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07669_ _03289_ _00121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06685__A1 _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_80_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09408_ ci_neuron.output_val_internal\[5\] _04633_ _04638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09339_ _04582_ _00507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09198__I _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08426__A2 _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07874__C ci_neuron.uut_simple_neuron.titan_id_5\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10114_ _00238_ net249 ci_neuron.uut_simple_neuron.titan_id_4\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10132__CLK net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10045_ _00530_ net169 ci_neuron.output_val_internal\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04923__B2 internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06979__A2 _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05020_ net37 _00706_ _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_113_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06971_ _02602_ _02604_ _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05922_ _01533_ _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09690_ _00277_ net222 ci_neuron.uut_simple_neuron.x3\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08710_ internal_ih.spi_rx_byte_i\[2\] _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05853_ _01456_ _01488_ _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08641_ _03915_ _04107_ _04113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_89_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05784_ _01444_ _01446_ _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08572_ _03950_ _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07523_ _03071_ _03134_ _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_49_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07454_ _03007_ _03009_ _03081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06405_ ci_neuron.uut_simple_neuron.x3\[9\] ci_neuron.uut_simple_neuron.x3\[10\]
+ _02050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07385_ _03012_ _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_79_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06336_ _01835_ _01952_ _01982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_79_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09124_ _04458_ _00416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06267_ _01915_ _00167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09055_ _04389_ _04400_ _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05218_ ci_neuron.uut_simple_neuron.x2\[9\] _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08006_ _03570_ _00148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06198_ _01847_ _01848_ _01849_ _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_12_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06198__A3 _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05149_ _00828_ _00224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09957_ _00472_ net76 ci_neuron.uut_simple_neuron.x0\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08908_ internal_ih.byte3\[7\] internal_ih.byte2\[7\] _04296_ _04298_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09392__I0 _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09888_ _00049_ net20 ci_neuron.value_i\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08839_ internal_ih.byte0\[1\] _04146_ _04258_ _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_68_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05881__A2 _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09391__I _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10028_ ci_neuron.input_memory\[1\]\[28\] net85 ci_neuron.uut_simple_neuron.titan_id_1\[30\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06897__A1 _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07170_ _02730_ _02800_ _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06121_ _01740_ _01776_ _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06052_ _01707_ _01708_ _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08470__I _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05003_ _00697_ _00049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09811_ _00390_ net53 internal_ih.byte7\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09742_ _00321_ net221 ci_neuron.uut_simple_neuron.x2\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06954_ _02576_ _02588_ _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06885_ _02518_ _02520_ _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_126_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09673_ _00260_ net261 ci_neuron.uut_simple_neuron.x3\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05905_ _01419_ _01420_ _01525_ _01564_ _01429_ _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_05836_ _01304_ _01355_ _01497_ _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08624_ _04055_ _04096_ _04097_ _04098_ _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_89_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05767_ _01328_ _01382_ _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08555_ _04040_ _02387_ _04028_ _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_25_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07506_ _03118_ _03132_ _03133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_85_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05560__A1 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05698_ _01218_ _01325_ _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08486_ _03957_ _03979_ _03981_ _00255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_53_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07437_ _02983_ _03062_ _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07368_ _02994_ _02971_ _02995_ _02996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06165__I ci_neuron.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06319_ _01903_ _01965_ _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_91_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09107_ ci_neuron.output_val_internal\[31\] ci_neuron.output_val_internal\[23\] ci_neuron.output_val_internal\[15\]
+ ci_neuron.output_val_internal\[7\] _04366_ _04367_ _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_103_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07299_ ci_neuron.uut_simple_neuron.x3\[23\] _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09038_ _04360_ _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08565__A1 _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09380__I3 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_110_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06670_ _02256_ _02299_ _02309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05621_ _01226_ ci_neuron.uut_simple_neuron.x2\[19\] _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_64_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05552_ _00886_ _01207_ _01219_ _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08340_ _03836_ _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05483_ _01133_ _01152_ _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08271_ _03790_ _03791_ _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_50_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07222_ _02821_ _02831_ _02851_ _02852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07153_ _02716_ _02782_ _02783_ _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_116_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06104_ _01756_ _01759_ _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07084_ _02712_ _02715_ _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06035_ _01657_ _01676_ _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout103 net104 net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08547__A1 _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout114 net116 net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout125 net127 net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout147 net164 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout136 net138 net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout158 net160 net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07986_ _03553_ _00145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout169 net171 net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06937_ _02570_ _02514_ _02571_ _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05781__A1 _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09725_ _00304_ net258 ci_neuron.uut_simple_neuron.x2\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09347__I0 _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09656_ _04827_ _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06868_ _02380_ _02503_ _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__05064__I _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08570__I1 _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08607_ _04019_ _04082_ _04083_ _04084_ _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_06799_ _02135_ _02394_ _02435_ _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_05819_ _01479_ _01480_ _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09587_ _00710_ _00713_ ci_neuron.interrupt_enabled _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08538_ _03943_ _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_92_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08469_ _03963_ _03964_ _03966_ _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_108_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06261__A2 _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09338__I0 _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08777__A1 _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06252__A2 _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07840_ _03430_ _00152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07771_ ci_neuron.uut_simple_neuron.titan_id_4\[22\] ci_neuron.uut_simple_neuron.titan_id_3\[22\]
+ _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06722_ _02321_ _02347_ _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09510_ _03848_ ci_neuron.input_memory\[1\]\[20\] ci_neuron.uut_simple_neuron.x2\[20\]
+ _02620_ _04716_ _04717_ _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_04983_ _00685_ _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07504__A2 _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06653_ _02289_ _02292_ _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_69_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09441_ ci_neuron.output_memory\[11\] _04650_ _04665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06584_ _02086_ _02189_ _02224_ _02225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_82_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05604_ _01263_ _01270_ _01271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09372_ _04606_ _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_35_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout33_I net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05535_ _01200_ _01203_ _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08323_ _03835_ _03836_ _03837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_62_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05466_ _01090_ _01094_ _01136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08254_ ci_neuron.uut_simple_neuron.x0\[9\] _03776_ _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__08923__I _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07205_ _02709_ _02760_ _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05397_ _01066_ _01023_ _01068_ _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08185_ _03717_ _03718_ _03719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07136_ _02639_ _02637_ _02765_ _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_113_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07067_ _02648_ _02699_ _02700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_30_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06018_ _01661_ _01675_ _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05059__I _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09568__I0 _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09193__A1 _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09708_ _00287_ net125 internal_ih.spi_rx_byte_i\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_07969_ ci_neuron.uut_simple_neuron.titan_id_2\[23\] ci_neuron.uut_simple_neuron.titan_id_5\[23\]
+ ci_neuron.uut_simple_neuron.titan_id_2\[22\] ci_neuron.uut_simple_neuron.titan_id_5\[22\]
+ _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09496__A2 _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09639_ ci_neuron.stream_o\[21\] ci_neuron.output_memory\[21\] _04816_ _04818_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_81_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_13_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08833__I _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06234__A2 _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10276_ _00569_ net133 ci_neuron.stream_o\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09681__CLK net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08782__I1 _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_100_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout168_I net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05320_ _00960_ _00990_ _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05251_ _00882_ _00902_ _00927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__04859__I0 internal_ih.byte4\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05182_ _00859_ _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06225__A2 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09990_ _00505_ net85 ci_neuron.input_memory\[1\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08941_ _04316_ _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08872_ _04277_ _00345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07823_ _03414_ _03416_ _03417_ _03418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07094__I _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07754_ ci_neuron.uut_simple_neuron.titan_id_4\[19\] ci_neuron.uut_simple_neuron.titan_id_3\[19\]
+ _03360_ _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_79_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04966_ _00676_ _00063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06705_ _02085_ _02343_ _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07685_ _03299_ _03300_ _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06636_ _02136_ _02233_ _02276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04897_ _00635_ _00019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09424_ ci_neuron.output_memory\[8\] _04650_ _04651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06567_ _02208_ _00232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09355_ _04591_ _00514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06498_ _02089_ _02095_ _02140_ _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_90_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05518_ _01096_ ci_neuron.uut_simple_neuron.x2\[16\] ci_neuron.uut_simple_neuron.x2\[17\]
+ _01187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_74_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09286_ _03974_ _04544_ _04552_ _00484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08306_ _03821_ _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05449_ _01119_ _01071_ _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08237_ _03741_ _03752_ _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_10_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08168_ _03692_ _03700_ _03703_ _03704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07119_ _02749_ _02750_ _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08099_ ci_neuron.uut_simple_neuron.titan_id_1\[15\] ci_neuron.uut_simple_neuron.titan_id_0\[15\]
+ _03647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10130_ _00200_ net265 ci_neuron.uut_simple_neuron.titan_id_3\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10061_ _00546_ net165 ci_neuron.output_val_internal\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05727__A1 _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08563__I _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07652__A1 ci_neuron.uut_simple_neuron.titan_id_4\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09547__I3 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10259_ _00552_ net151 ci_neuron.stream_o\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout285_I net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07470_ _02725_ _03096_ _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06421_ _02065_ _00229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06352_ _01964_ _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09140_ _04466_ _00424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_118_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06283_ _01874_ _01904_ _01930_ _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05303_ ci_neuron.uut_simple_neuron.x2\[11\] _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09071_ _04377_ _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08022_ ci_neuron.uut_simple_neuron.titan_id_1\[3\] ci_neuron.uut_simple_neuron.titan_id_0\[3\]
+ _03582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05234_ ci_neuron.uut_simple_neuron.x2\[10\] _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05165_ _00834_ _00843_ _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05096_ _00777_ _00200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09973_ _00488_ net178 ci_neuron.input_memory\[1\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_90_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08924_ internal_ih.byte4\[6\] internal_ih.byte3\[6\] _04306_ _04307_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08855_ _04267_ _00338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_129_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07806_ _03397_ _03399_ _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08786_ _04017_ _00977_ _04225_ _04228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07737_ _03342_ _03343_ _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05998_ _01527_ _01626_ _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04949_ internal_ih.byte0\[1\] _00665_ _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_95_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07668_ _03287_ _03288_ _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06685__A2 _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07599_ _02604_ _02630_ _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06619_ _01836_ _02212_ _02259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09407_ _04630_ _04636_ _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_109_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09338_ _04104_ ci_neuron.input_memory\[1\]\[27\] _04578_ _04582_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09269_ _04139_ _04535_ spi_interface_cvonk.state\[2\] _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10113_ _00237_ net243 ci_neuron.uut_simple_neuron.titan_id_4\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10044_ _00529_ net170 ci_neuron.output_val_internal\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_102_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07625__A1 _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_113_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06970_ _02125_ _02127_ _02603_ _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_05921_ _01574_ _01578_ _01580_ _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05852_ _01460_ _01487_ _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08640_ _04112_ _00278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05783_ _01400_ _01404_ _01445_ _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08571_ _04054_ _00267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07522_ _03073_ _03147_ _03148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07453_ _03011_ _03015_ _03079_ _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06404_ _01961_ _02002_ _02048_ _02049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_76_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07384_ _02936_ _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09123_ ci_neuron.uut_simple_neuron.titan_id_6\[5\] _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07616__A1 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06335_ _01976_ _01978_ _01981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_79_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06266_ _01912_ _01914_ _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09054_ ci_neuron.output_val_internal\[26\] ci_neuron.output_val_internal\[18\] ci_neuron.output_val_internal\[10\]
+ ci_neuron.output_val_internal\[2\] _04390_ _04391_ _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_44_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05217_ _00869_ _00893_ _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08005_ ci_neuron.uut_simple_neuron.titan_id_2\[29\] ci_neuron.uut_simple_neuron.titan_id_5\[29\]
+ _03569_ _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06197_ _01837_ _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05148_ _00806_ _00827_ _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05067__I _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05079_ _00759_ _00761_ _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09956_ _00471_ net86 ci_neuron.uut_simple_neuron.x0\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08907_ _04297_ _00360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09887_ _00048_ net19 ci_neuron.value_i\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09392__I1 ci_neuron.input_memory\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08838_ _04257_ _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09541__A1 ci_neuron.output_memory\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08769_ _03974_ _04209_ _04217_ _00302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_28_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05094__A1 _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07457__I ci_neuron.uut_simple_neuron.x3\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput5 net5 spi_poci_o vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_31_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10027_ ci_neuron.input_memory\[1\]\[27\] net85 ci_neuron.uut_simple_neuron.titan_id_1\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06897__A2 _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout248_I net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06120_ _01743_ _01775_ _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06051_ _01618_ _01620_ _01671_ _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_30_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05002_ internal_ih.byte3\[0\] _00696_ _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_74_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08949__I1 internal_ih.byte5\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09810_ _00389_ net54 internal_ih.byte7\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06953_ _02587_ _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09741_ _00320_ net223 ci_neuron.uut_simple_neuron.x2\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_129_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05904_ _01427_ _01525_ _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06884_ _02464_ _02462_ _02519_ _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_126_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05615__I _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09672_ _00259_ net261 ci_neuron.uut_simple_neuron.x3\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05835_ _01400_ _01444_ _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08623_ ci_neuron.value_i\[26\] _03965_ _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05766_ _01423_ _01419_ _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_49_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08554_ _03996_ _04037_ _04038_ _04039_ _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_25_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07505_ _03120_ _03131_ _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_85_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05697_ _01254_ _01325_ _01360_ _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08485_ _01900_ _03980_ _03981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07436_ _02991_ _02988_ _03063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07367_ _02922_ _02961_ _02995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06318_ _01960_ _01964_ _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09106_ _04417_ ci_neuron.stream_o\[7\] ci_neuron.stream_o\[23\] _04418_ _04446_
+ _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_07298_ _02731_ _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09037_ _04359_ _04384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06249_ _01830_ _01881_ _01897_ _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_60_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09939_ _00454_ net176 ci_neuron.uut_simple_neuron.x0\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08836__I _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09373__S0 _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05620_ _01261_ _01272_ _01285_ _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07650__I _03274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07819__A1 ci_neuron.uut_simple_neuron.titan_id_4\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05551_ _01105_ _01151_ _01192_ _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_59_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05482_ _01148_ _01151_ _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_58_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08270_ _03782_ _03784_ _03786_ _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_50_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07221_ _02794_ _02820_ _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08619__I0 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07152_ _02718_ _02759_ _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06103_ _01669_ _01757_ _01758_ _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07083_ _01835_ _01871_ _02714_ _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06034_ _01689_ _01690_ _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout104 net106 net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09595__I1 ci_neuron.output_memory\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout115 net116 net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout126 net127 net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout137 net138 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout148 net150 net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout159 net160 net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07985_ _03551_ _03552_ _03553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06936_ _02474_ _02513_ _02571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05345__I _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09724_ _00303_ net257 ci_neuron.uut_simple_neuron.x2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_2_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06867_ _02500_ _02502_ _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_87_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09655_ ci_neuron.stream_o\[28\] ci_neuron.output_memory\[28\] _04826_ _04827_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05818_ _01433_ _01291_ _01380_ _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_69_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08606_ ci_neuron.value_i\[23\] _04013_ _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06798_ _02096_ _02279_ _02435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_38_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09586_ _04787_ _00549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05749_ _01255_ _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08537_ _03797_ _03798_ _04015_ _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08468_ ci_neuron.value_i\[3\] _03965_ _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07419_ _01867_ _01936_ _03045_ _03046_ _03047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_80_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08399_ ci_neuron.uut_simple_neuron.x0\[28\] _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09283__I0 _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_107_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07277__A2 _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05288__A1 _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09397__I _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06788__A1 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07770_ _03373_ _00109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04982_ _00599_ _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06721_ _02315_ _02316_ _02317_ _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_91_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09440_ _04649_ _04661_ _04663_ _04664_ _00526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06652_ _02291_ _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_69_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06583_ _02222_ _02223_ _02224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_87_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05603_ _00741_ _01265_ _01269_ _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09371_ _03935_ _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_35_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05534_ _01201_ _01202_ _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_86_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08322_ ci_neuron.uut_simple_neuron.x0\[19\] _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout26_I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08253_ ci_neuron.uut_simple_neuron.x0\[10\] _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_15_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07204_ _02781_ _02834_ _02835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_117_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05465_ _01090_ _01094_ _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05396_ _01067_ _01024_ _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08184_ ci_neuron.uut_simple_neuron.titan_id_1\[30\] ci_neuron.uut_simple_neuron.titan_id_0\[30\]
+ _03718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07135_ _02700_ _02705_ _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07066_ _02649_ _02698_ _02699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06017_ _01674_ _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09568__I1 ci_neuron.input_memory\[1\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09193__A2 _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05203__A1 _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07968_ _03531_ _03536_ _03538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06919_ _02445_ _02501_ _02553_ _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09707_ _00286_ net131 internal_ih.spi_rx_byte_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_97_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07899_ _03477_ _03479_ _03480_ _03481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__06703__A1 _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09638_ _04817_ _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09569_ _04768_ _04774_ _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08456__A1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09256__I0 _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10275_ _00568_ net142 ci_neuron.stream_o\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05250_ _00922_ _00925_ _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__04859__I1 internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05181_ _00858_ _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08940_ internal_ih.byte5\[5\] internal_ih.byte4\[5\] _04312_ _04316_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_110_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08871_ internal_ih.byte1\[7\] internal_ih.byte0\[7\] _04275_ _04277_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07822_ ci_neuron.uut_simple_neuron.titan_id_4\[30\] ci_neuron.uut_simple_neuron.titan_id_3\[30\]
+ _03417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07753_ _03350_ _03355_ _03356_ _03358_ _03359_ _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_04965_ internal_ih.byte1\[0\] _00675_ _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06704_ _02051_ _02186_ _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_07684_ ci_neuron.uut_simple_neuron.titan_id_4\[7\] ci_neuron.uut_simple_neuron.titan_id_3\[7\]
+ _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04896_ internal_ih.byte4\[4\] _00633_ _00634_ internal_ih.byte0\[4\] _00635_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06635_ _01898_ _02274_ _02275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_94_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09423_ _04599_ _04650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09354_ _04589_ _04590_ _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06566_ _02166_ _02167_ _02207_ _02208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08305_ ci_neuron.uut_simple_neuron.x0\[16\] _03821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06497_ _02090_ _02139_ _02140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05517_ _01185_ _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09285_ ci_neuron.input_memory\[1\]\[4\] _04549_ _04552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05448_ _01065_ _01069_ _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08236_ _03748_ _03749_ _03760_ _03747_ _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_10_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08167_ ci_neuron.uut_simple_neuron.titan_id_1\[27\] ci_neuron.uut_simple_neuron.titan_id_0\[27\]
+ _03702_ _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07118_ _01863_ _02665_ _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05379_ _01049_ _01050_ _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_42_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07413__A2 _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05424__A1 _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08098_ _03646_ _00070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07049_ _02555_ _02681_ _02682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10060_ _00545_ net103 ci_neuron.output_val_internal\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07101__A1 _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08601__A1 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10258_ _00551_ net151 ci_neuron.stream_o\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05718__A2 _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10189_ _00087_ net44 ci_neuron.uut_simple_neuron.titan_id_2\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout180_I net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06420_ _02027_ _02026_ _02064_ _02065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_69_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06351_ _01896_ _01967_ _01996_ _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_71_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06282_ _01878_ _01903_ _01930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_84_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05302_ ci_neuron.uut_simple_neuron.x2\[6\] _00861_ _00975_ _00976_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_72_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09483__I3 _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09070_ _04378_ _04413_ _04414_ _00406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05233_ _00863_ _00892_ _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08021_ _03581_ _00077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05164_ _00821_ _00842_ _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_77_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout6 net7 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05406__A1 _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05095_ _00772_ _00776_ _00777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09972_ _00487_ net178 ci_neuron.input_memory\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08923_ _04290_ _04306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08854_ internal_ih.byte1\[0\] internal_ih.byte0\[0\] _04264_ _04267_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07805_ _03402_ _00115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05997_ _01611_ _01625_ _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08785_ _04010_ _04211_ _04227_ _00308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07736_ ci_neuron.uut_simple_neuron.titan_id_4\[16\] ci_neuron.uut_simple_neuron.titan_id_3\[16\]
+ _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04948_ _00666_ _00033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07331__A1 _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07667_ ci_neuron.uut_simple_neuron.titan_id_4\[5\] ci_neuron.uut_simple_neuron.titan_id_3\[5\]
+ _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04879_ internal_ih.byte4\[7\] internal_ih.byte3\[7\] _00601_ _00623_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06618_ _02256_ _02257_ _02258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07598_ _02178_ _03219_ _03222_ _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09406_ _03742_ ci_neuron.input_memory\[1\]\[5\] _00795_ _01900_ _04622_ _04623_
+ _04636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_48_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06549_ _02184_ _02190_ _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09337_ _04581_ _00506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09268_ _04138_ _04140_ _04540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_23_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07634__A2 _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08219_ _03746_ _00195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09199_ _03742_ _04500_ _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10112_ _00236_ net287 ci_neuron.uut_simple_neuron.titan_id_4\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10043_ _00528_ net166 ci_neuron.output_val_internal\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07570__A1 _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07322__A1 _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05920_ _01472_ _01532_ _01579_ _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05851_ _01450_ _01490_ _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08570_ _04052_ _02445_ _04053_ _04054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07521_ _03133_ _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05782_ _01396_ _01399_ _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07452_ _03016_ _03020_ _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08484__I _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07864__A2 ci_neuron.uut_simple_neuron.titan_id_5\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07383_ _02859_ _03010_ _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06403_ _01964_ _02001_ _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06334_ _01980_ _00169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09122_ _04457_ _00415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08813__A1 _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06265_ _01886_ _01913_ _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_72_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09053_ _04383_ ci_neuron.stream_o\[2\] ci_neuron.stream_o\[18\] _04384_ _04398_
+ _04399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_115_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06196_ _01822_ _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_05216_ ci_neuron.uut_simple_neuron.x2\[0\] _00838_ _00892_ _00893_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08004_ _03565_ _03567_ _03568_ _03569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05147_ _00824_ _00826_ _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05078_ _00760_ _00757_ _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09955_ _00470_ net88 ci_neuron.uut_simple_neuron.x0\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08906_ internal_ih.byte3\[6\] internal_ih.byte2\[6\] _04296_ _04297_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09886_ _00047_ net22 ci_neuron.value_i\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09392__I2 _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08837_ _04256_ _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07552__A1 _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08768_ _00768_ _04214_ _04217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_28_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07719_ _03331_ _00099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08699_ internal_ih.spi_tx_byte_o\[5\] _04136_ _04157_ internal_ih.spi_rx_byte_i\[5\]
+ _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_0_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07855__A2 ci_neuron.uut_simple_neuron.titan_id_5\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05094__A2 _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08569__I _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10026_ ci_neuron.input_memory\[1\]\[26\] net76 ci_neuron.uut_simple_neuron.titan_id_1\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06346__A2 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07543__A1 ci_neuron.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09296__A1 _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06050_ _00936_ _01706_ _01668_ _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_2_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05001_ _00685_ _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06952_ _02583_ _02586_ _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09740_ _00319_ net223 ci_neuron.uut_simple_neuron.x2\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
.ends

