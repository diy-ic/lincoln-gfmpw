* NGSPICE file created from titan.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

.subckt titan spi_clock_i spi_cs_i spi_pico_i spi_poci_o sys_clock_i vdd vss
X_05903_ _01561_ _01562_ _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06883_ _02418_ _02461_ _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09671_ _00258_ clknet_leaf_51_sys_clock_i ci_neuron.uut_simple_neuron.x3\[8\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05834_ _01162_ _01200_ _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08622_ _03889_ _03879_ _04081_ _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05765_ _01427_ _01428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08553_ ci_neuron.value_i\[15\] _04001_ _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07504_ _03123_ _03130_ _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08484_ _03968_ _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07435_ _02979_ _03060_ _03062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05696_ _01252_ _01324_ _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_65_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07366_ _02962_ _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_128_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07297_ _02873_ _02877_ _02925_ _02926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06317_ ci_neuron.uut_simple_neuron.x3\[8\] _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_98_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09105_ _04360_ _04445_ _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06248_ _01877_ _01896_ _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_103_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05076__A2 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09036_ _04361_ _04383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06179_ _01827_ _01830_ _01831_ _01832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09211__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold340 internal_ih.byte7\[7\] net373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold362 _04588_ net395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold351 internal_ih.byte7\[5\] net384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold373 ci_neuron.uut_simple_neuron.x0\[17\] net406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold384 ci_neuron.uut_simple_neuron.x0\[29\] net417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold395 internal_ih.byte4\[4\] net428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09938_ _00453_ clknet_leaf_73_sys_clock_i ci_neuron.uut_simple_neuron.x0\[9\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_5_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09869_ _00060_ net26 ci_neuron.value_i\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_107_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09373__S1 _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrebuffer7 _02311_ net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_106_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09202__A1 _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_69_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10009_ net58 clknet_leaf_81_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05550_ _00859_ _01178_ _01174_ _01218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_82_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05481_ _01097_ _01150_ _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07220_ _02789_ _02848_ _02849_ _02850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08619__I1 _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07151_ _02718_ _02759_ _02782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06102_ _00747_ ci_neuron.uut_simple_neuron.x2\[29\] _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09441__A1 ci_neuron.output_memory\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07082_ _01835_ _02713_ _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06033_ _01650_ _01679_ _01690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_93_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold472_I internal_ih.byte0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07984_ ci_neuron.uut_simple_neuron.titan_id_2\[26\] net695 _03552_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06935_ _02472_ _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08555__I0 _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09723_ _00302_ clknet_leaf_67_sys_clock_i ci_neuron.uut_simple_neuron.x2\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06866_ _02388_ _02501_ _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_hold737_I internal_ih.byte0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09654_ _04810_ _04826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_96_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05817_ _01327_ _01478_ _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08605_ _03864_ _04077_ _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06797_ _02376_ _02432_ _02433_ _02434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09585_ _04607_ net229 _04785_ _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_120_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05748_ _01361_ _01409_ _01410_ _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08536_ _04024_ _00262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05679_ _01342_ _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08467_ _03950_ _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08483__A2 _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07418_ _01988_ _01991_ _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08398_ _03902_ _00188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07349_ _02977_ _02974_ _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_135_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09019_ internal_ih.data_pointer\[1\] _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_131_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08621__B _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold170 ci_neuron.stream_o\[26\] net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold192 ci_neuron.output_val_internal\[25\] net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold181 _00517_ net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__04980__A1 internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09510__I2 ci_neuron.uut_simple_neuron.x2\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06237__A1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06788__A2 _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07737__A1 _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05212__A2 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04981_ _00684_ _00039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06720_ _02358_ _00235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08757__I _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04971__A1 internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06651_ _02044_ _02290_ _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_78_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05602_ _00937_ _01266_ _01268_ _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06582_ _02188_ _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05181__I _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09370_ _04604_ _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_129_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05533_ _01123_ _01162_ _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08321_ net617 _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05464_ _01131_ _01107_ _01133_ _01056_ _01134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_75_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08252_ _03775_ _00199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07203_ _02784_ _02833_ _02834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_132_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05395_ _00934_ _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_104_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08183_ _03692_ _03700_ _03712_ _03716_ _03717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_07134_ _02647_ _02765_ _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07065_ _02652_ _02697_ _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_101_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06016_ _01665_ _01673_ _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07728__A1 ci_neuron.uut_simple_neuron.titan_id_4\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09568__I2 _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07967_ net461 _00142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_113_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06918_ _02498_ _02552_ _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08528__I0 _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09706_ net119 clknet_leaf_103_sys_clock_i internal_ih.spi_rx_byte_i\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_07898_ ci_neuron.uut_simple_neuron.titan_id_2\[11\] ci_neuron.uut_simple_neuron.titan_id_5\[11\]
+ _03480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04962__A1 internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06703__A2 _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06849_ _02440_ _02456_ _02485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09637_ ci_neuron.stream_o\[20\] net323 _04816_ _04817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_104_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09568_ _03915_ ci_neuron.input_memory\[1\]\[29\] _01751_ ci_neuron.uut_simple_neuron.x3\[29\]
+ _04760_ _04761_ _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_08519_ ci_neuron.value_i\[10\] _03971_ _04009_ _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_33_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09499_ ci_neuron.output_memory\[19\] _04698_ _04715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_137_Right_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_135_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_122_Left_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09405__A1 ci_neuron.output_memory\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06219__A1 _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10274_ _00567_ clknet_leaf_108_sys_clock_i ci_neuron.stream_o\[16\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_131_Left_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_140_Left_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05180_ net33 _00837_ _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_77_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08870_ _04276_ _00344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07821_ ci_neuron.uut_simple_neuron.titan_id_4\[30\] ci_neuron.uut_simple_neuron.titan_id_3\[30\]
+ _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07752_ ci_neuron.uut_simple_neuron.titan_id_4\[18\] ci_neuron.uut_simple_neuron.titan_id_3\[18\]
+ _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04964_ _00664_ _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06703_ _02332_ _02341_ _02342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07683_ net523 _00123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_88_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08686__A2 _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04895_ _00627_ _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06634_ _01907_ _02273_ _02274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06697__A1 _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09422_ _04597_ _04649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09353_ net730 _04352_ _04590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06565_ _02203_ _02206_ _02207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06449__A1 _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08304_ _03820_ _00176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06496_ _02094_ _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05516_ _01096_ _01149_ _01184_ _01185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09284_ _04551_ _00483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05447_ _01116_ _01117_ _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08235_ _03752_ ci_neuron.uut_simple_neuron.x0\[7\] _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_31_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05378_ _01012_ _01020_ _00961_ _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08166_ _03696_ _03701_ _03702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07117_ _02175_ _02193_ _02749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08097_ _03643_ _03645_ _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07048_ ci_neuron.uut_simple_neuron.x3\[21\] ci_neuron.uut_simple_neuron.x3\[22\]
+ _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_11_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08999_ net283 _04341_ _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_48_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08921__I0 internal_ih.byte4\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_95_sys_clock_i clknet_4_10_0_sys_clock_i clknet_leaf_95_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_124_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08601__A2 _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10257_ _00000_ clknet_leaf_127_sys_clock_i ci_neuron.stream_enabled vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10188_ _00086_ clknet_leaf_4_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[30\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06350_ _01994_ _01995_ _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_57_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06281_ _01928_ _01929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05301_ ci_neuron.uut_simple_neuron.x2\[7\] ci_neuron.uut_simple_neuron.x2\[8\] _00975_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05232_ _00894_ _00897_ _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08770__I _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08020_ net606 ci_neuron.uut_simple_neuron.titan_id_0\[3\] _03580_ _03581_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_25_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold703 _03434_ net736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05163_ _00840_ _00841_ _00842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold736 _01900_ net769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold714 ci_neuron.uut_simple_neuron.titan_id_2\[15\] net747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold725 _01751_ net758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout7 net8 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold747 ci_neuron.uut_simple_neuron.titan_id_4\[25\] net780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_05094_ _00736_ _00774_ _00775_ _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09971_ _00486_ clknet_leaf_67_sys_clock_i ci_neuron.input_memory\[1\]\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold758 ci_neuron.uut_simple_neuron.titan_id_0\[28\] net791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold769 ci_neuron.uut_simple_neuron.titan_id_5\[30\] net802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08922_ net463 _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08853_ net382 _00337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_137_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07804_ net601 _03401_ _03402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05996_ _01609_ _01627_ _01653_ _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08784_ _00911_ _04221_ _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04917__B2 internal_ih.byte1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_139_sys_clock_i_I clknet_4_0_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07735_ net694 _00102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04947_ internal_ih.byte0\[0\] _00665_ _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07666_ _03283_ _03285_ _03286_ _03287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_79_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_04878_ _00622_ _00031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_36_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09405_ ci_neuron.output_memory\[5\] _04628_ _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07597_ _03220_ _03221_ _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06617_ _02245_ _02202_ _02244_ _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
Xclkbuf_leaf_137_sys_clock_i clknet_4_0_0_sys_clock_i clknet_leaf_137_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_118_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06548_ _02086_ _02189_ _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09336_ _04099_ net92 _04578_ _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07095__A1 _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09267_ _04537_ _04139_ _04538_ _04535_ _04539_ _00478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_06479_ _00163_ _02121_ _02122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08218_ _03740_ _03742_ _03745_ _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_117_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09198_ _04499_ _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08149_ _03684_ _03686_ _03687_ _03688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10111_ _00235_ clknet_leaf_44_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_112_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10042_ net104 clknet_leaf_112_sys_clock_i ci_neuron.output_val_internal\[11\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_145_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold41 ci_neuron.input_memory\[1\]\[13\] net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_54_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold30 net650 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_145_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold63 net821 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold52 ci_neuron.input_memory\[1\]\[4\] net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold74 ci_neuron.output_val_internal\[8\] net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold96 ci_neuron.uut_simple_neuron.titan_id_6\[12\] net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold85 _04154_ net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07322__A2 _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_44_sys_clock_i clknet_4_7_0_sys_clock_i clknet_leaf_44_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_85_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08822__A2 _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09622__I1 ci_neuron.output_memory\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_58_sys_clock_i_I clknet_4_15_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05850_ _01453_ _01489_ _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09550__A3 _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer17 _02287_ net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05454__I _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07520_ _03135_ _03139_ _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05781_ _01236_ _01408_ _01443_ _01444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
Xrebuffer28 _02003_ net448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_85_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08510__A1 ci_neuron.value_i\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07451_ _03076_ _03026_ _03077_ _03078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06402_ _01926_ _02004_ _02046_ _02047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07382_ _03009_ _03007_ _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_9_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06333_ _01943_ _01979_ _01980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09121_ net208 _04457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06264_ _01884_ _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_89_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09052_ _04385_ _04397_ _04398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold500 _03361_ net533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06195_ _01825_ _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_103_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05215_ _00891_ _00892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold511 _03833_ net544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_4_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_127_sys_clock_i_I clknet_4_2_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08003_ net773 net554 _03568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold544 _03370_ net577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_130_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05146_ _00802_ _00825_ _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold522 spi_interface_cvonk.SS_r\[0\] net666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__09613__I1 ci_neuron.output_memory\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold533 ci_neuron.uut_simple_neuron.titan_id_0\[31\] net566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold577 ci_neuron.uut_simple_neuron.titan_id_3\[23\] net610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_111_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold566 _03314_ net599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold555 _03652_ net588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold588 _03807_ net621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold599 ci_neuron.uut_simple_neuron.titan_id_4\[8\] net632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05077_ _00753_ _00760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09954_ _00469_ clknet_leaf_14_sys_clock_i ci_neuron.uut_simple_neuron.x0\[25\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08905_ _04290_ _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09885_ _00046_ net22 ci_neuron.value_i\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08836_ _04185_ _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_127_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09392__I3 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05979_ _01593_ _01596_ _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08767_ _04216_ _00301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07718_ net456 ci_neuron.uut_simple_neuron.titan_id_3\[13\] _03330_ _03331_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08698_ _04133_ net201 _04161_ _00287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07649_ _03225_ _03270_ _03273_ _03274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_79_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09319_ _04571_ _00498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08804__A2 _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06291__A2 _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09604__I1 net316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10025_ net88 clknet_leaf_31_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08786__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05554__A1 _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06833__I _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05000_ _00695_ _00048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10007__D net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06951_ _02301_ _02307_ _02585_ _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_94_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05902_ _01538_ _01542_ _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09670_ _00257_ clknet_leaf_51_sys_clock_i ci_neuron.uut_simple_neuron.x3\[7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06882_ _02515_ _02517_ _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08621_ _03879_ _04082_ _03890_ _04096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05833_ _01493_ _01494_ _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05545__A1 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05764_ _01419_ _01420_ _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08552_ _03817_ _04030_ _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_clkbuf_leaf_115_sys_clock_i_I clknet_4_9_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07503_ _00162_ _03129_ _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08483_ ci_neuron.value_i\[5\] _03952_ _03978_ _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_9_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07434_ _03061_ _00246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_122_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05695_ _01323_ _01348_ _01349_ _01284_ _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_07365_ _02963_ _02970_ _02992_ _02993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_116_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07296_ _02862_ _02872_ _02925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06316_ _01900_ _01932_ _01962_ _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_98_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09104_ _04419_ ci_neuron.stream_o\[15\] _04445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06247_ net36 _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09035_ _04355_ _04382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06178_ _01826_ _01828_ _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold341 _04338_ net374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold352 _04336_ net385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold330 _04791_ net363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_99_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05129_ _00773_ _00795_ _00767_ _00809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
Xhold374 _03832_ net407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold396 net744 net429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold363 ci_neuron.uut_simple_neuron.x0\[26\] net396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold385 _03912_ net418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09937_ _00452_ clknet_leaf_73_sys_clock_i ci_neuron.uut_simple_neuron.x0\[8\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07525__A2 _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09868_ _00059_ net25 ci_neuron.value_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09514__A3 _04726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08819_ _04094_ _01573_ _04246_ _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09799_ _00378_ clknet_leaf_144_sys_clock_i internal_ih.byte6\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09278__A2 _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07289__A1 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_15_0_sys_clock_i clknet_0_sys_clock_i clknet_4_15_0_sys_clock_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_134_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer8 _01108_ net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05775__A1 _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08713__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09505__A3 _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10008_ net59 clknet_leaf_62_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_69_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05480_ _01149_ _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_67_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_17_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07150_ _02780_ _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_89_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07081_ _01936_ _01868_ _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_112_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06101_ _00738_ _01751_ _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_81_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06032_ _01654_ _01678_ _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_103_sys_clock_i_I clknet_4_8_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09722_ _00301_ clknet_leaf_66_sys_clock_i ci_neuron.uut_simple_neuron.x2\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07983_ net790 _03548_ _03550_ _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06934_ _02526_ _02568_ _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06865_ ci_neuron.uut_simple_neuron.x3\[18\] ci_neuron.uut_simple_neuron.x3\[19\]
+ _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_2_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09653_ _04825_ _00578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05816_ ci_neuron.uut_simple_neuron.x2\[23\] _01380_ _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08604_ _04081_ _04082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09584_ _04786_ _00548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06796_ _02378_ _02397_ _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08535_ _04023_ _02226_ _03969_ _04024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05747_ _01366_ _01393_ _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05678_ _01342_ _01328_ _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_65_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08466_ _03730_ _03958_ _03953_ _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_9_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_35_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07417_ _01988_ _01958_ _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_92_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08397_ _03898_ _03901_ _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_21_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07348_ _02847_ _02975_ _02976_ _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07443__A1 _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07279_ _02897_ _02908_ _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_135_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09018_ internal_ih.data_pointer\[0\] _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07994__A2 ci_neuron.uut_simple_neuron.titan_id_5\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09196__A1 _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold171 _04403_ net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold160 _00520_ net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_44_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_130_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold182 ci_neuron.stream_o\[27\] net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold193 _00541_ net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_73_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06182__A1 ci_neuron.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10110__D _00234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09510__I3 _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_22_sys_clock_i_I clknet_4_6_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04980_ internal_ih.byte1\[7\] _00680_ _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06650_ net448 _02141_ _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_05601_ _01267_ _01265_ _01268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_8_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08974__S _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06581_ _02186_ _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05532_ _01158_ _01161_ _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08320_ net544 _03834_ _00178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05463_ _01058_ _01132_ _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08251_ _03770_ _03772_ _03774_ _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07202_ _02789_ _02792_ _02832_ _02833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_117_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05394_ _00999_ _01066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08182_ _03715_ _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07133_ _02699_ _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07425__A1 _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07064_ _02656_ _02696_ _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07976__A2 net823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06015_ _01616_ _01672_ _01673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09568__I3 ci_neuron.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07966_ net460 _03536_ _03537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06917_ _02551_ _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08528__I1 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09705_ net162 clknet_leaf_103_sys_clock_i internal_ih.spi_rx_byte_i\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07897_ ci_neuron.uut_simple_neuron.titan_id_2\[11\] ci_neuron.uut_simple_neuron.titan_id_5\[11\]
+ _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09636_ _04810_ _04816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06848_ _02476_ _02483_ _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06779_ _02361_ _02400_ _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_104_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09567_ net196 _04766_ _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08518_ _03945_ _04008_ _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09498_ _04697_ _04711_ _04713_ _04714_ _00534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xclkbuf_leaf_94_sys_clock_i clknet_4_10_0_sys_clock_i clknet_leaf_94_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_137_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08449_ _03941_ _03947_ _03949_ _00250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07299__I ci_neuron.uut_simple_neuron.x3\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06219__A2 _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_115_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10273_ _00566_ clknet_leaf_99_sys_clock_i ci_neuron.stream_o\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_10_sys_clock_i_I clknet_4_4_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09495__I2 _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07407__A1 _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_5_sys_clock_i_I clknet_4_1_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06630__A2 _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07820_ net741 _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07751_ _03342_ _03343_ _03357_ _03358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06702_ _02223_ _02340_ _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_04963_ _00674_ _00062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06288__I _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07682_ _03299_ net522 _03301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_88_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04894_ _00605_ _00633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06633_ _01994_ _02236_ _02272_ _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_94_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_136_sys_clock_i clknet_4_2_0_sys_clock_i clknet_leaf_136_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09421_ _04627_ _04643_ _04647_ _04648_ _00523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06564_ _02204_ _02205_ _02206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09352_ _00583_ _04353_ _04589_ _00513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05515_ ci_neuron.uut_simple_neuron.x2\[17\] _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08303_ _03814_ _03819_ _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06495_ _01995_ _02097_ _02137_ _02138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09283_ _03967_ net56 _04543_ _04551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_119_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05446_ _01074_ _01077_ _01115_ _01117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_90_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08234_ _03759_ _00197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_31_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05377_ _01012_ _01020_ _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08165_ ci_neuron.uut_simple_neuron.titan_id_1\[27\] ci_neuron.uut_simple_neuron.titan_id_0\[27\]
+ _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_132_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07116_ _02743_ _02747_ _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08096_ net547 _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07047_ _02551_ _02624_ _02679_ _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_100_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08998_ _04348_ _00400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07949_ _03520_ _03521_ _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_43_sys_clock_i clknet_4_7_0_sys_clock_i clknet_leaf_43_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09619_ net342 _00563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_39_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07637__A1 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10256_ _00550_ clknet_leaf_127_sys_clock_i ci_neuron.interrupt_enabled vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10187_ _00085_ clknet_leaf_3_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09078__B1 ci_neuron.stream_o\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06280_ _01853_ _01906_ _01927_ _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05300_ _00973_ _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_86_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05231_ _00889_ _00899_ _00906_ _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05162_ _00813_ _00817_ _00839_ _00841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
Xhold726 _00910_ net759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold715 _03494_ net748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold737 internal_ih.byte0\[5\] net808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_12_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout8 net16 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold704 _03436_ net737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold748 _03388_ net781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_122_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05093_ _00744_ _00758_ _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09970_ _00485_ clknet_leaf_74_sys_clock_i ci_neuron.input_memory\[1\]\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold759 ci_neuron.uut_simple_neuron.titan_id_0\[25\] net792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08921_ internal_ih.byte4\[5\] net462 _04301_ _04305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08852_ internal_ih.byte0\[7\] net381 _04264_ _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07803_ _03396_ _03397_ _03400_ _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05995_ _01568_ _01629_ _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08783_ _04226_ _00307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07734_ _03342_ _03343_ _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04946_ _00664_ _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07665_ ci_neuron.uut_simple_neuron.titan_id_4\[4\] ci_neuron.uut_simple_neuron.titan_id_3\[4\]
+ _03286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06616_ _02241_ _02243_ _02256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_95_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_9_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_04877_ internal_ih.byte7\[6\] _00616_ _00621_ _00597_ _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_36_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09404_ _04627_ _04629_ _04632_ _04634_ _00520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_07596_ _03152_ _03211_ _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06547_ _02186_ _02188_ _02189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09335_ _04580_ _00505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06478_ _02079_ _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09266_ net249 _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_132_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05429_ _00969_ _01005_ _01052_ _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_08217_ _03743_ _03744_ _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09197_ _04486_ _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08148_ net719 net796 _03687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08079_ _03627_ _03628_ _03629_ _03630_ _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_30_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10110_ _00234_ clknet_leaf_42_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_112_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10041_ net114 clknet_leaf_112_sys_clock_i ci_neuron.output_val_internal\[10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_145_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold31 net668 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_145_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold64 net820 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold42 net761 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold53 net806 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold86 _00285_ net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold97 internal_ih.spi_tx_byte_o\[6\] net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold75 _00524_ net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_85_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05097__A1 _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09910__CLK net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06340__B _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _00135_ clknet_leaf_117_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xrebuffer18 _02688_ net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05780_ _01411_ _01442_ _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_89_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer29 _02871_ net499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_1
XFILLER_0_107_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08510__A2 _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07450_ _03004_ _03021_ _03077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06401_ _02044_ _02045_ _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07381_ _02868_ _03008_ _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08649__I0 _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06332_ _01976_ _01978_ _01979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_84_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08781__I _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09120_ _04456_ _00414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09051_ _04358_ ci_neuron.stream_o\[10\] _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06263_ _01890_ _01909_ _01911_ _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08002_ net773 net554 _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06194_ _01820_ _01845_ _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_05214_ _00811_ _00846_ ci_neuron.uut_simple_neuron.x2\[8\] _00891_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xhold501 internal_ih.spi_rx_byte_i\[5\] net534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_142_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05145_ _00782_ _00819_ _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold545 net822 net578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold512 _00178_ net545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold523 spi_interface_cvonk.MOSI_r\[0\] net668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_40_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold534 ci_neuron.uut_simple_neuron.titan_id_2\[1\] net567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold578 _03379_ net611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold567 ci_neuron.uut_simple_neuron.titan_id_4\[28\] net600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06588__A1 _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold556 _03655_ net589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_60_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05076_ _00737_ _00745_ _00759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09953_ _00468_ clknet_leaf_12_sys_clock_i ci_neuron.uut_simple_neuron.x0\[24\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold589 ci_neuron.uut_simple_neuron.titan_id_1\[4\] net622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_hold662_I ci_neuron.uut_simple_neuron.titan_id_5\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08904_ net360 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09884_ _00045_ net19 ci_neuron.value_i\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08835_ _04255_ _00330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_127_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10203__D _00099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08766_ _03967_ _00758_ _04208_ _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05978_ _01634_ _01636_ _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07717_ _03326_ _03327_ _03329_ _03330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09385__S0 _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08697_ internal_ih.spi_rx_byte_i\[5\] _04148_ _04161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04929_ internal_ih.byte6\[1\] _00652_ _00653_ internal_ih.byte2\[1\] _00655_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07648_ _03271_ _03214_ _03272_ _03213_ _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_0_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07579_ _02079_ _03204_ _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09318_ _04059_ net89 _04567_ _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06815__A2 _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09249_ _04528_ _00471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10024_ net91 clknet_leaf_11_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[26\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06751__A1 ci_neuron.uut_simple_neuron.x3\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05242__A1 _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06950_ _02578_ _02584_ _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06881_ _02422_ _02460_ _02516_ _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05901_ _01523_ _01537_ _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input3_I spi_pico_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05832_ _01448_ _01451_ _01491_ _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08620_ _04095_ _00275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05763_ _01421_ _01424_ _01386_ _01425_ _01343_ _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_08551_ _03809_ _04036_ _03825_ _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07502_ _03126_ _03128_ _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05694_ _01358_ _00212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08482_ _03965_ _03976_ _03977_ _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08495__A1 _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07433_ _02990_ _03060_ _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_122_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_4_0_sys_clock_i clknet_0_sys_clock_i clknet_4_4_0_sys_clock_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07364_ _02966_ _02969_ _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_99_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout8_I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09103_ _04415_ net236 _04444_ _00409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07295_ _02879_ _02883_ _02923_ _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06315_ _01959_ _01961_ _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_98_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06246_ _01894_ _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09034_ _04370_ _04381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold320 internal_ih.byte7\[6\] net353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_130_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06177_ _01829_ _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold342 ci_neuron.input_memory\[1\]\[31\] net375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold353 ci_neuron.uut_simple_neuron.x0\[12\] net386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold331 ci_neuron.stream_o\[15\] net364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05128_ _00787_ _00807_ _00808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold375 ci_neuron.uut_simple_neuron.titan_id_3\[1\] net408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold364 internal_ih.byte7\[3\] net397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold386 internal_ih.byte3\[4\] net419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05059_ _00743_ _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09936_ _00451_ clknet_leaf_76_sys_clock_i ci_neuron.uut_simple_neuron.x0\[7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold397 internal_ih.byte6\[5\] net430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_51_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09867_ _00058_ net25 ci_neuron.value_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06733__A1 _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07590__I _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08818_ _04224_ _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09798_ _00377_ clknet_leaf_143_sys_clock_i internal_ih.byte5\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08749_ _04194_ net290 _00296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_138_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08635__B _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09310__I _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer9 net55 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05285__I _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10007_ net61 clknet_leaf_82_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_69_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08477__A1 _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07080_ _02710_ _02711_ _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06100_ _01755_ _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_124_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06031_ _01648_ _01681_ _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05463__A1 _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07982_ _03545_ _03550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06933_ _02567_ _02528_ _02568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__06963__A1 _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09721_ _00300_ clknet_leaf_67_sys_clock_i ci_neuron.uut_simple_neuron.x2\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06864_ _02383_ _02448_ _02499_ _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_2_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold458_I internal_ih.byte4\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09652_ net215 net315 _04821_ _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06795_ _02378_ _02397_ _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05815_ _01474_ _01476_ _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08603_ _03863_ _04077_ _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09583_ _04605_ net350 _04785_ _04786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_2_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05746_ _01366_ _01393_ _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08468__A1 ci_neuron.value_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08534_ _04020_ _04022_ _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_49_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_93_sys_clock_i clknet_4_11_0_sys_clock_i clknet_leaf_93_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05677_ ci_neuron.uut_simple_neuron.x2\[21\] _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08465_ _03729_ _03958_ _03963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_07416_ _03042_ _03043_ _03044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08396_ _03895_ _03899_ _03900_ _03894_ _03901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_21_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07347_ _02850_ _02909_ _02976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07278_ _02899_ _02907_ _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_135_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09017_ _04355_ _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06229_ _01873_ _01878_ _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold150 spi_interface_cvonk.buffer\[7\] net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold161 ci_neuron.uut_simple_neuron.titan_id_6\[0\] net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold194 internal_ih.spi_rx_byte_i\[2\] net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold183 _04413_ net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold172 ci_neuron.uut_simple_neuron.titan_id_6\[11\] net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09919_ _00016_ net6 ci_neuron.address_i\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_29_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08631__A1 _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09187__A2 _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07198__A1 _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05600_ _01226_ _01264_ _01267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_135_sys_clock_i clknet_4_2_0_sys_clock_i clknet_leaf_135_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_145_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06580_ _02191_ _02194_ _02220_ _02221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_87_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05531_ _01166_ _01199_ _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_24_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05462_ _01106_ _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08250_ _03773_ _03766_ _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07201_ _02821_ _02831_ _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08181_ _03707_ _03713_ _03712_ _03703_ _03714_ _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_6_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07132_ _02763_ _02761_ _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_132_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05393_ _00932_ _01064_ _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_sys_clock_i_I sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07063_ _02658_ _02695_ _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_42_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06014_ _01666_ _01671_ _01672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07965_ ci_neuron.uut_simple_neuron.titan_id_2\[23\] ci_neuron.uut_simple_neuron.titan_id_5\[23\]
+ _03536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06916_ ci_neuron.uut_simple_neuron.x3\[19\] _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09704_ _00283_ clknet_leaf_103_sys_clock_i internal_ih.spi_rx_byte_i\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_42_sys_clock_i clknet_4_7_0_sys_clock_i clknet_leaf_42_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_97_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07896_ net729 _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09635_ net368 _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06847_ _02479_ _02482_ _02483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06778_ _02415_ _00236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_104_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09566_ _04765_ _04767_ _04770_ _04772_ _00544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05729_ _01388_ _01392_ _01393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08517_ _04006_ _04007_ _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09497_ net120 _04705_ _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_137_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08448_ _02898_ _03948_ _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08379_ _03882_ _03876_ _03885_ _03881_ _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_18_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10272_ _00565_ clknet_leaf_111_sys_clock_i ci_neuron.stream_o\[14\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09495__I3 _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07407__A2 _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_95_sys_clock_i_I clknet_4_10_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07750_ ci_neuron.uut_simple_neuron.titan_id_4\[16\] ci_neuron.uut_simple_neuron.titan_id_3\[16\]
+ _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06394__A2 _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04962_ internal_ih.byte0\[7\] _00670_ _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06701_ _02337_ _02339_ _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_07681_ net521 ci_neuron.uut_simple_neuron.titan_id_3\[7\] _03300_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04893_ _00632_ _00018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06632_ _01995_ _02135_ _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_88_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09420_ net168 _04633_ _04648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06563_ _02160_ _02158_ _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09351_ _04145_ _04152_ _04352_ _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_118_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05514_ _01175_ _01182_ _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09282_ _03961_ _04544_ _04550_ _00482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08302_ _03816_ _03818_ _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07646__A2 _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06494_ _02135_ _02136_ _02137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08233_ _03754_ _03756_ _03758_ _03759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA_fanout24_I net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05445_ _01074_ _01077_ _01115_ _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_90_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05376_ _00860_ _01044_ _01047_ _01048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08164_ _03693_ _03698_ _03700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09643__I0 ci_neuron.stream_o\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07115_ _02225_ _02746_ _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08095_ ci_neuron.uut_simple_neuron.titan_id_1\[15\] net546 _03644_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07046_ _02555_ _02623_ _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_30_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08997_ net282 _04341_ _04348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07948_ _03517_ _03518_ _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07879_ ci_neuron.uut_simple_neuron.titan_id_2\[8\] net304 _03461_ _03462_ _03464_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_48_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09618_ net341 ci_neuron.output_memory\[12\] _04805_ _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_39_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09549_ net219 _04749_ _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10255_ _00549_ clknet_leaf_120_sys_clock_i ci_neuron.normalised_stream_write_address\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10186_ _00084_ clknet_leaf_3_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07325__A1 _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07013__I _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_83_sys_clock_i_I clknet_4_14_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_62_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05230_ _00890_ _00898_ _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_126_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05161_ _00813_ _00817_ _00839_ _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_80_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold727 ci_neuron.uut_simple_neuron.x2\[23\] net760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_80_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold705 ci_neuron.uut_simple_neuron.x2\[22\] net738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold716 ci_neuron.uut_simple_neuron.x0\[5\] net749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout9 net10 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold749 ci_neuron.uut_simple_neuron.titan_id_4\[27\] net782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05092_ _00773_ _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold738 _02928_ net771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08920_ net420 _00366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_71_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08851_ net465 _00336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07802_ ci_neuron.uut_simple_neuron.titan_id_4\[27\] ci_neuron.uut_simple_neuron.titan_id_3\[27\]
+ _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05994_ _01649_ _01651_ _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08782_ _04003_ _00896_ _04225_ _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07733_ net693 net580 _03343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04945_ _00599_ _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07664_ ci_neuron.uut_simple_neuron.titan_id_4\[4\] ci_neuron.uut_simple_neuron.titan_id_3\[4\]
+ _03285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07867__A2 ci_neuron.uut_simple_neuron.titan_id_5\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04876_ internal_ih.byte4\[6\] internal_ih.byte3\[6\] _00601_ _00621_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06615_ _02247_ _02255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09403_ net192 _04633_ _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07595_ _03155_ _03210_ _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06546_ _02094_ _02187_ _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_80_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08816__A1 _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09334_ _04094_ net88 _04578_ _04580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06477_ _02113_ _02063_ _02112_ _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_118_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09265_ _04166_ _04138_ _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05428_ _00939_ _01054_ _01091_ _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_62_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08216_ _03733_ _03737_ _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09196_ _03974_ _04494_ _04498_ _00448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05359_ _01004_ _01022_ _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08147_ net719 net796 _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_141_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08078_ ci_neuron.uut_simple_neuron.titan_id_1\[11\] ci_neuron.uut_simple_neuron.titan_id_0\[11\]
+ _03630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07029_ _02178_ _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_112_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10040_ net112 clknet_leaf_112_sys_clock_i ci_neuron.output_val_internal\[9\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_145_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold32 net665 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_145_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold43 ci_neuron.input_memory\[1\]\[10\] net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold54 net793 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold65 net700 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07307__A1 _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold98 _04164_ net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold87 ci_neuron.output_val_internal\[18\] net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold76 ci_neuron.output_val_internal\[15\] net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_119_Left_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_14_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09480__A1 ci_neuron.output_memory\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05097__A2 _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_128_Left_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10238_ _00134_ clknet_leaf_117_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10169_ _00095_ clknet_leaf_84_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_71_sys_clock_i_I clknet_4_12_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_137_Left_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xrebuffer19 _02612_ net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09223__I _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06400_ _02003_ _02045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07380_ ci_neuron.uut_simple_neuron.x3\[26\] ci_neuron.uut_simple_neuron.x3\[27\]
+ _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06331_ _01890_ _01944_ _01917_ _01977_ _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_44_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06262_ _01827_ _01884_ _01910_ _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09050_ _04378_ net191 _04396_ _00404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05213_ _00742_ _00862_ _00870_ _00890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_5_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08001_ _03566_ _00147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06193_ _01842_ _01844_ _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xhold502 ci_neuron.uut_simple_neuron.titan_id_1\[27\] net535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_4_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold524 ci_neuron.uut_simple_neuron.titan_id_3\[15\] net557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_102_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05144_ _00810_ _00823_ _00824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold513 ci_neuron.uut_simple_neuron.titan_id_0\[15\] net546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__09885__CLK net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold568 _03399_ net601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold579 _03383_ net612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06588__A2 _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05075_ _00757_ _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold557 ci_neuron.uut_simple_neuron.titan_id_5\[4\] net590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold546 _03787_ net579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09952_ _00467_ clknet_4_4_0_sys_clock_i ci_neuron.uut_simple_neuron.x0\[23\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_140_sys_clock_i_I clknet_4_0_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08903_ internal_ih.byte3\[5\] net359 _04291_ _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07537__A1 _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09883_ _00043_ net21 ci_neuron.value_i\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08834_ net505 _04143_ _04254_ _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_127_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08765_ _03961_ _04209_ _04215_ _00300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05977_ _01076_ _01592_ _01635_ _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07716_ ci_neuron.uut_simple_neuron.titan_id_4\[12\] ci_neuron.uut_simple_neuron.titan_id_3\[12\]
+ _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_140_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09385__S1 _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08696_ net200 _04136_ _04157_ internal_ih.spi_rx_byte_i\[4\] _04160_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_04928_ _00654_ _00008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07647_ _03146_ _03143_ _03272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04859_ internal_ih.byte4\[1\] internal_ih.byte3\[1\] _00608_ _00609_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07578_ _02088_ _02103_ _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_0_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06529_ _02130_ _02151_ _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09317_ _04570_ _00497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09248_ _04104_ _03892_ _04525_ _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09179_ _04485_ _04206_ _04486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09517__A2 _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10023_ net81 clknet_leaf_11_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09043__I internal_ih.data_pointer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09453__A1 ci_neuron.output_memory\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09205__A1 _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06880_ _02424_ _02459_ _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05900_ _01389_ _01558_ _01559_ _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05831_ _01492_ _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05762_ _00749_ _01384_ _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08550_ _04030_ _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07501_ _02074_ _03127_ _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05693_ _01355_ _01357_ _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08481_ _03739_ _03963_ _03741_ _03977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_92_sys_clock_i clknet_4_11_0_sys_clock_i clknet_leaf_92_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07432_ _03059_ _02991_ _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_122_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08792__I _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_18_sys_clock_i_I clknet_4_3_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07363_ _02974_ _02977_ _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09102_ net130 _04427_ _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07294_ _02856_ _02853_ _02878_ _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06314_ _01960_ _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_98_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06245_ _01891_ _01893_ _01894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09033_ net207 _04378_ _04380_ _00403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_142_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06176_ _01819_ _01828_ _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__05481__A2 _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold310 internal_ih.byte7\[0\] net343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_130_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05127_ _00792_ _00797_ _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold343 ci_neuron.uut_simple_neuron.titan_id_5\[12\] net376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold321 _04337_ net354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold332 _04809_ net365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold376 _03420_ net409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold354 ci_neuron.uut_simple_neuron.x0\[24\] net387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold387 _04304_ net420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold365 _04334_ net398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05058_ _00742_ _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09935_ _00450_ clknet_leaf_76_sys_clock_i ci_neuron.uut_simple_neuron.x0\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold398 internal_ih.byte4\[6\] net431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09866_ _00055_ net25 ci_neuron.value_i\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08817_ net739 _04236_ _04245_ _00322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08183__A1 _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09797_ _00376_ clknet_leaf_143_sys_clock_i internal_ih.byte5\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08748_ net289 _04202_ _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_107_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08486__A2 _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08679_ net68 _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_83_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08797__I0 _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08877__I _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10006_ net60 clknet_leaf_82_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06724__A2 _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07921__A1 _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_134_sys_clock_i clknet_4_2_0_sys_clock_i clknet_leaf_134_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_114_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09501__I _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_132_Right_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06030_ _01652_ _01680_ _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08788__I0 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07981_ _03549_ _00144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06932_ _02538_ _02540_ _02566_ _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_09720_ _00299_ clknet_leaf_31_sys_clock_i ci_neuron.uut_simple_neuron.x2\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04974__A1 internal_ih.byte1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold186_I ci_neuron.output_val_internal\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41_sys_clock_i clknet_4_7_0_sys_clock_i clknet_leaf_41_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06863_ _02388_ _02498_ _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_2_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09651_ _04824_ _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06794_ _02365_ _02430_ _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05814_ _00748_ _01475_ _01476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08602_ _03986_ _04079_ _04080_ _00272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09582_ _04599_ _00730_ _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05745_ _01406_ _01407_ _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08533_ _03789_ _04006_ _04021_ _03959_ _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__06479__A1 _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08468__A2 _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05676_ _01338_ _01340_ _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08464_ _03957_ _03961_ _03962_ _00252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07415_ _02953_ _02959_ _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08395_ net396 _03891_ _03900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_9_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07346_ _02850_ _02909_ _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_102_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07277_ _02902_ _02906_ _02907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_135_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09016_ _04358_ ci_neuron.stream_o\[0\] ci_neuron.stream_o\[16\] _04359_ _04363_
+ _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_33_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06228_ ci_neuron.uut_simple_neuron.x3\[5\] _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06159_ ci_neuron.uut_simple_neuron.x2\[31\] _01812_ _01813_ _01814_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xhold162 ci_neuron.uut_simple_neuron.x0\[8\] net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold140 ci_neuron.uut_simple_neuron.x0\[4\] net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold151 _04169_ net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold195 _00332_ net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold184 _00406_ net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold173 ci_neuron.stream_o\[24\] net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09918_ _00015_ net19 ci_neuron.address_i\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08156__A1 _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09849_ _00428_ clknet_leaf_115_sys_clock_i ci_neuron.output_memory\[17\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08631__A2 _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04956__A1 internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05920__A3 _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05530_ _01124_ _01198_ _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05461_ _01088_ _01095_ _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07200_ _02824_ _02830_ _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05392_ _01032_ _01063_ _01064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08180_ net799 ci_neuron.uut_simple_neuron.titan_id_0\[29\] _03714_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07131_ _02649_ _02698_ _02762_ _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08083__B1 _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07062_ _02694_ _02668_ _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_11_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06013_ _00936_ _01668_ _01670_ _01671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04947__A1 internal_ih.byte0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold470_I internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07964_ net459 _03534_ _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06915_ _02380_ _02503_ _02549_ _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07895_ ci_neuron.uut_simple_neuron.titan_id_2\[11\] net728 _03477_ _03478_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09703_ net255 clknet_leaf_132_sys_clock_i net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06846_ _01824_ _02481_ _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_hold735_I _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09634_ ci_neuron.stream_o\[19\] net367 _04811_ _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06777_ _02410_ _02414_ _02415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_104_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05372__A1 _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08466__B _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09565_ ci_neuron.output_val_internal\[28\] _04771_ _04772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05728_ _01389_ _01391_ _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08516_ _03782_ _03997_ _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09496_ _04701_ _04712_ _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_136_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05659_ _01146_ _01223_ _01287_ _01324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_08447_ _03940_ _03948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_137_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08378_ _03874_ _03875_ _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07329_ _01968_ _02957_ _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09661__I1 net361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10271_ _00564_ clknet_leaf_111_sys_clock_i ci_neuron.stream_o\[13\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_100_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09252__S _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05363__A1 _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05418__A2 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_90_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06918__A2 _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04929__B2 internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04961_ _00673_ _00061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06700_ _02283_ _02338_ _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07680_ _03295_ _03297_ _03298_ _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_04892_ internal_ih.byte4\[3\] _00625_ _00628_ internal_ih.byte0\[3\] _00632_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06631_ _02219_ _02269_ _02270_ _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_88_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06562_ _02154_ _02157_ _02204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09350_ net395 _00512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05513_ _01179_ _01181_ _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08301_ _03811_ _03817_ _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09281_ net90 _04549_ _04550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06493_ _02096_ _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08232_ _03742_ _03754_ _03757_ _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05444_ _01078_ _01114_ _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05375_ _01017_ _01046_ _01047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08163_ _03699_ _00083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_132_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07114_ _02234_ _02745_ _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08094_ _03639_ _03640_ _03642_ _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_70_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07045_ _02495_ _02626_ _02677_ _02678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_63_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08996_ _04347_ _00399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07582__A2 _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07947_ ci_neuron.uut_simple_neuron.titan_id_2\[20\] net483 _03520_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08906__I0 internal_ih.byte3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07878_ net565 _00157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08531__A1 ci_neuron.value_i\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06829_ _02463_ _02465_ _02466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_97_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09617_ _04789_ _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_39_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09548_ _04746_ _04756_ _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09479_ _04674_ _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06845__A1 _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09011__A2 internal_ih.data_pointer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10254_ _00548_ clknet_leaf_120_sys_clock_i ci_neuron.normalised_stream_write_address\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10185_ _00083_ clknet_leaf_14_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07325__A2 _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08522__A1 _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05336__A1 _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05749__I _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05160_ _00733_ _00835_ _00838_ _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08589__A1 _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold706 _01473_ net739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold728 ci_neuron.input_memory\[1\]\[24\] net805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold717 ci_neuron.input_memory\[1\]\[1\] net795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_110_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05091_ _00760_ _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold739 ci_neuron.uut_simple_neuron.titan_id_1\[31\] net772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09002__A2 _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08850_ internal_ih.byte0\[6\] net464 _04264_ _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07801_ net600 ci_neuron.uut_simple_neuron.titan_id_3\[28\] _03399_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08761__A1 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05993_ _01650_ _01631_ _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08781_ _04224_ _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07732_ _03338_ _03340_ _03341_ _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_04944_ _00663_ _00016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05327__A1 _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07663_ net636 _00120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04875_ _00620_ _00030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06614_ _02254_ _00233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_36_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09402_ _04610_ _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07594_ _02808_ _03217_ _03218_ _03219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_88_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09333_ _04579_ _00504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06545_ ci_neuron.uut_simple_neuron.x3\[12\] ci_neuron.uut_simple_neuron.x3\[13\]
+ _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08816__A2 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06476_ _02070_ _02116_ _02118_ _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09264_ net249 _04127_ _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05427_ _01097_ _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08215_ _03730_ _03740_ _03743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09195_ _03740_ _04491_ _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08146_ net720 _00080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05358_ _01004_ _01022_ _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07252__A1 _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05289_ ci_neuron.uut_simple_neuron.x2\[9\] _00910_ ci_neuron.uut_simple_neuron.x2\[11\]
+ _00963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_08077_ ci_neuron.uut_simple_neuron.titan_id_1\[11\] ci_neuron.uut_simple_neuron.titan_id_0\[11\]
+ ci_neuron.uut_simple_neuron.titan_id_1\[10\] ci_neuron.uut_simple_neuron.titan_id_0\[10\]
+ _03629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_15_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07028_ _01846_ _02659_ _02660_ _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_112_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_145_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold55 net775 net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold44 net757 net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_54_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold33 net686 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08979_ net354 _00392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09741__D _00320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold99 _00289_ net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold88 _00534_ net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold66 net831 net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold77 _00531_ net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_97_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09304__I0 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06953__I _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10237_ _00133_ clknet_leaf_92_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10168_ _00094_ clknet_leaf_84_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10099_ _00165_ clknet_leaf_55_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_91_sys_clock_i clknet_4_11_0_sys_clock_i clknet_leaf_91_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_107_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06330_ _01940_ _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06261_ _01871_ _01883_ _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05212_ _00835_ _00888_ _00869_ _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_4_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08000_ net773 net554 _03565_ _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_143_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06192_ ci_neuron.uut_simple_neuron.x3\[1\] _01843_ _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05143_ _00818_ _00819_ _00822_ _00784_ _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
Xhold525 _03339_ net558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold514 _03644_ net547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold503 _03698_ net536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold536 _03423_ net569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold547 ci_neuron.uut_simple_neuron.titan_id_3\[16\] net580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold569 _03402_ net602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_96_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05074_ _00756_ _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09951_ _00466_ clknet_leaf_18_sys_clock_i ci_neuron.uut_simple_neuron.x0\[22\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold558 _03437_ net591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08982__A1 _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08902_ net335 _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07537__A2 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09882_ _00042_ net19 ci_neuron.value_i\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05548__A1 _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08833_ _04192_ _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_127_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05976_ _01556_ _01591_ _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08764_ _00774_ _04214_ _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07715_ net679 _00098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04927_ internal_ih.byte6\[0\] _00652_ _00653_ internal_ih.byte2\[0\] _00654_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_140_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08695_ _04134_ net239 _04159_ _00286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07646_ _03141_ _03066_ _03271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_94_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04858_ _00600_ _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_137_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07577_ _03201_ _03202_ _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06528_ _02168_ _02169_ _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09316_ _04052_ net71 _04567_ _04570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09247_ _04527_ _00470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09462__A2 _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06459_ _02102_ _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09178_ _03934_ _03936_ _04485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08129_ _03668_ _03669_ _03671_ _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_102_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_56_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10022_ net67 clknet_leaf_12_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_133_sys_clock_i clknet_4_2_0_sys_clock_i clknet_leaf_133_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_40_sys_clock_i clknet_4_5_0_sys_clock_i clknet_leaf_40_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05830_ _01448_ _01451_ _01491_ _01492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07500_ _02081_ _02480_ _03127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05761_ _01105_ _01422_ _01371_ _01373_ _01423_ _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05692_ _01304_ _01314_ _01356_ _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08480_ _03739_ _03741_ _03963_ _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_49_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07431_ _02993_ _03055_ _03058_ _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_122_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07362_ _02988_ _02989_ _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06313_ ci_neuron.uut_simple_neuron.x3\[7\] _01960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_84_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09101_ net235 _04416_ _04442_ _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07293_ _02885_ _02895_ _02921_ _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_98_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06244_ _01892_ _01841_ _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09032_ net125 _04379_ _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07207__A1 _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06175_ ci_neuron.uut_simple_neuron.x3\[1\] ci_neuron.uut_simple_neuron.x3\[2\] _01828_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_5_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold311 _04330_ net344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold300 _04808_ net333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05126_ _00804_ _00805_ _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold344 _03482_ net377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold333 ci_neuron.uut_simple_neuron.x0\[11\] net366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold322 ci_neuron.stream_o\[10\] net355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold366 net750 net399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold355 _03874_ net388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold377 internal_ih.byte4\[7\] net410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_05057_ _00741_ _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09934_ _00449_ clknet_leaf_76_sys_clock_i ci_neuron.uut_simple_neuron.x0\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold388 internal_ih.byte5\[5\] net421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold399 internal_ih.byte2\[2\] net432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08707__A1 _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09865_ _00044_ net27 ci_neuron.value_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08816_ _04089_ _04237_ _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_59_sys_clock_i clknet_4_14_0_sys_clock_i clknet_leaf_59_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_51_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09796_ _00375_ clknet_leaf_142_sys_clock_i internal_ih.byte5\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05959_ _01472_ _01532_ _01579_ _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08747_ _04193_ net210 _04202_ _00295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_107_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08678_ _04145_ _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07629_ _03252_ _03253_ _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06497__A2 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08797__I1 _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10005_ net57 clknet_leaf_81_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_69_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09875__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07988__A2 net695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07980_ _03546_ _03548_ _03549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06931_ _02544_ _02565_ _02566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09650_ net203 net328 _04821_ _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_124_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06862_ ci_neuron.uut_simple_neuron.x3\[18\] _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08601_ _02805_ _04011_ _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06793_ _02427_ _02429_ _02430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05813_ ci_neuron.uut_simple_neuron.x2\[24\] _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09581_ _04765_ _04781_ _04783_ _04784_ _00547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05744_ _00934_ _01395_ _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08532_ _03799_ _04006_ _04021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06479__A2 _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08463_ _01849_ _03948_ _03962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07414_ _02956_ _02958_ _03042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05675_ _01186_ _01287_ _01339_ _01146_ _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07212__I _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08394_ _03889_ _03891_ _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07345_ _02973_ _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_116_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07276_ _02904_ _02905_ _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06227_ _01876_ _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09015_ _04360_ _04362_ _04363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06158_ _01464_ _01462_ _01454_ _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold130 net818 net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold141 _03739_ net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold152 _00290_ net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_06089_ _01700_ _01719_ _01745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05109_ _00780_ _00782_ _00783_ _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold185 ci_neuron.uut_simple_neuron.titan_id_6\[18\] net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold174 _04372_ net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold163 ci_neuron.output_memory\[29\] net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold196 ci_neuron.normalised_stream_write_address\[1\] net229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09917_ _00014_ net6 ci_neuron.address_i\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09848_ _00427_ clknet_leaf_115_sys_clock_i ci_neuron.output_memory\[16\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05914__A1 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09779_ _00358_ clknet_leaf_1_sys_clock_i internal_ih.byte3\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09512__I _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05460_ _01129_ _01095_ _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05391_ _01034_ _01038_ _01062_ _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_83_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07130_ _02652_ _02697_ _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04892__A1 internal_ih.byte4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07061_ _02693_ _02671_ _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_101_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06012_ _00738_ _01669_ _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07963_ _03530_ _03531_ _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06914_ _02547_ _02548_ _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07894_ _03473_ _03474_ _03476_ _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09702_ net64 clknet_leaf_101_sys_clock_i internal_ih.spi_rx_byte_i\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06845_ _02038_ _02480_ _02481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09633_ net262 _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09564_ _04704_ _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06776_ _02308_ _02412_ _02413_ _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_104_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08515_ _04005_ _03998_ _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09422__I _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05727_ _00864_ _01207_ _01390_ _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_77_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09495_ _03841_ ci_neuron.input_memory\[1\]\[18\] _01227_ _02616_ _04691_ _04692_
+ _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA_clkbuf_leaf_79_sys_clock_i_I clknet_4_14_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05658_ _01321_ _01295_ _01322_ _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_93_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08446_ ci_neuron.value_i\[0\] _03944_ _03946_ _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_137_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08377_ _03884_ _00185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07328_ _02374_ _02395_ _02957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05589_ _01255_ _01220_ _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_73_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07259_ _02282_ _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_103_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10270_ _00563_ clknet_leaf_98_sys_clock_i ci_neuron.stream_o\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09913__CLK net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08860__I0 net481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08612__S _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05100__I net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09565__A1 ci_neuron.output_val_internal\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09507__I _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04960_ internal_ih.byte0\[6\] _00670_ _00673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06630_ _02221_ _02239_ _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04891_ _00631_ _00017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_88_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06561_ _02199_ _02202_ _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06303__A1 _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06492_ _02093_ _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05512_ _01147_ _01180_ _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09280_ _04545_ _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08300_ _03808_ _03810_ _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05443_ _01081_ _01113_ _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08231_ _03748_ _03749_ _03747_ _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_4_11_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06854__A2 _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold211_I ci_neuron.output_val_internal\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05374_ _00982_ _01045_ _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08162_ _03697_ net536 _03699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_31_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07113_ _02379_ _02685_ _02744_ _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08093_ ci_neuron.uut_simple_neuron.titan_id_1\[14\] ci_neuron.uut_simple_neuron.titan_id_0\[14\]
+ _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_70_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07044_ _02622_ _02676_ _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_31_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09417__I _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07031__A2 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_67_sys_clock_i_I clknet_4_12_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08995_ net281 _04340_ _04347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07946_ net485 _00139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07877_ _03461_ _03462_ _03463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08531__A2 _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06828_ _02408_ _02405_ _02464_ _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_143_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09616_ net326 _00562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_39_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06759_ _02393_ _02396_ _02397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09547_ _03890_ ci_neuron.input_memory\[1\]\[26\] _01579_ _03083_ _04738_ _04739_
+ _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_39_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09478_ _04696_ _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08429_ ci_neuron.address_i\[0\] _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_136_sys_clock_i_I clknet_4_2_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10253_ _00151_ clknet_leaf_4_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10184_ _00082_ clknet_leaf_14_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[26\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_90_sys_clock_i clknet_4_11_0_sys_clock_i clknet_leaf_90_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08522__A2 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08286__A1 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08589__A2 _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold707 ci_neuron.uut_simple_neuron.titan_id_4\[30\] net740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold718 _01839_ net751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_25_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05090_ _00763_ _00771_ _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold729 _01264_ net762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_122_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04870__I1 internal_ih.byte3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07800_ _03398_ _00114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08780_ _04207_ _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_127_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05992_ _01604_ _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07731_ ci_neuron.uut_simple_neuron.titan_id_4\[15\] net557 _03341_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04943_ internal_ih.byte6\[7\] _00658_ _00659_ internal_ih.byte2\[7\] _00663_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07662_ net635 ci_neuron.uut_simple_neuron.titan_id_3\[4\] _03283_ _03284_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_04874_ internal_ih.byte7\[5\] _00616_ _00619_ _00597_ _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06613_ _02250_ _02253_ _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07593_ _02933_ _03012_ _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09401_ _04630_ _04631_ _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06544_ _02091_ _02143_ _02185_ _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09332_ _04089_ net91 _04578_ _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_145_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06475_ _02072_ _02115_ _02118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_leaf_55_sys_clock_i_I clknet_4_15_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09263_ _04127_ _04535_ _04536_ _00477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05426_ _01096_ _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08214_ _03741_ _03742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09194_ _03734_ _04489_ _04497_ _00447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05357_ _00996_ _01025_ _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08145_ net719 ci_neuron.uut_simple_neuron.titan_id_0\[24\] _03684_ _03685_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_15_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07252__A2 _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05288_ _00961_ _00892_ _00942_ _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__05263__A1 _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08076_ _03619_ _03624_ _03628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07027_ _02128_ _02603_ _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_112_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold23 net555 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05015__A1 internal_ih.byte3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10233__D _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold56 net794 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold45 net774 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold34 net568 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_54_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_132_sys_clock_i clknet_4_2_0_sys_clock_i clknet_leaf_132_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08978_ net353 internal_ih.byte6\[6\] _04257_ _04337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07929_ _03498_ _03503_ _03505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold89 ci_neuron.output_memory\[3\] net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold78 ci_neuron.output_val_internal\[9\] net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold67 ci_neuron.uut_simple_neuron.titan_id_6\[24\] net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_124_sys_clock_i_I clknet_4_3_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06190__B _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05585__I _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10236_ _00132_ clknet_leaf_86_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_5_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10167_ _00093_ clknet_leaf_84_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08896__I _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10098_ _00164_ clknet_leaf_63_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06809__A2 _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06260_ _01895_ _01899_ _01908_ _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_127_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05493__A1 _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05211_ _00887_ _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06191_ ci_neuron.uut_simple_neuron.x3\[2\] _01838_ _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__08806__I0 _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08580__B _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05142_ _00821_ _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold515 _03646_ net548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold526 ci_neuron.uut_simple_neuron.titan_id_0\[12\] net559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold504 spi_interface_cvonk.SCLK_r\[0\] net650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold548 _03345_ net581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_122_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold537 ci_neuron.uut_simple_neuron.titan_id_5\[19\] net570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05073_ ci_neuron.uut_simple_neuron.x2\[3\] _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09950_ _00465_ clknet_leaf_18_sys_clock_i ci_neuron.uut_simple_neuron.x0\[21\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold559 _03439_ net592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08982__A2 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08901_ internal_ih.byte3\[4\] net334 _04291_ _04294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_58_sys_clock_i clknet_4_15_0_sys_clock_i clknet_leaf_58_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09881_ _00041_ net22 ci_neuron.value_i\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08832_ _04253_ _00329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_43_sys_clock_i_I clknet_4_7_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05975_ _01449_ _01633_ _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08763_ _04210_ _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07714_ _03326_ net678 _03328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08498__A1 _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04926_ _00626_ _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08694_ internal_ih.spi_rx_byte_i\[4\] _04149_ _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_140_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07645_ _03239_ _03260_ _03269_ _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_04857_ _00607_ _00025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07576_ _02074_ _03127_ _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06527_ _01831_ _02129_ _02169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09315_ _04569_ _00496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06458_ _02101_ _02100_ _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09246_ _04099_ _03890_ _04525_ _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05409_ _01038_ _01062_ _01080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06389_ _01993_ _02011_ _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09177_ _00587_ _04187_ _04189_ _04353_ _00443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08128_ ci_neuron.uut_simple_neuron.titan_id_1\[20\] ci_neuron.uut_simple_neuron.titan_id_0\[20\]
+ _03671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08059_ net563 _00093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_56_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10021_ net75 clknet_leaf_12_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_112_sys_clock_i_I clknet_4_10_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09340__I _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05475__A1 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10219_ _00116_ clknet_leaf_3_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05760_ _01375_ _01337_ _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05691_ _01300_ _01303_ _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_12_0_sys_clock_i clknet_0_sys_clock_i clknet_4_12_0_sys_clock_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_59_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07430_ _02918_ _03056_ _03057_ _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_122_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07361_ _02979_ _02984_ _02989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06312_ _01903_ _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_84_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09100_ _04356_ _04439_ _04441_ _04411_ _04442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07292_ _02855_ _02884_ _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07455__A2 _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09031_ _04377_ _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06243_ _01820_ _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_98_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_31_sys_clock_i_I clknet_4_5_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_131_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06174_ _01826_ _01827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_68_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold301 internal_ih.byte2\[4\] net334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_05125_ _00778_ _00800_ _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold312 internal_ih.byte5\[7\] net345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA_hold493_I internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold323 _04803_ net356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold334 ci_neuron.output_memory\[19\] net367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold378 ci_neuron.uut_simple_neuron.titan_id_4\[9\] net411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold345 _03483_ net378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold356 _03876_ net389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold367 internal_ih.byte7\[4\] net400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05056_ _00740_ _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09933_ _00448_ clknet_leaf_79_sys_clock_i ci_neuron.uut_simple_neuron.x0\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold389 _04316_ net422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09864_ _00033_ net25 ci_neuron.value_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08815_ _04244_ _00321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_51_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09425__I _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09795_ _00374_ clknet_leaf_141_sys_clock_i internal_ih.byte5\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05958_ ci_neuron.uut_simple_neuron.x2\[1\] _01581_ _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_77_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08746_ internal_ih.received_byte_count\[5\] net209 _04199_ _04202_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_36_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05889_ _01547_ _01549_ _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_107_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08677_ net515 _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04909_ internal_ih.byte5\[1\] _00640_ _00641_ internal_ih.byte1\[1\] _00643_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_4_9_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07628_ _03194_ _03209_ _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09677__CLK clknet_4_13_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07559_ _02504_ _03101_ _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_100_sys_clock_i_I clknet_4_8_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_86_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09229_ _04517_ _00462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08504__I _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_95_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10004_ net85 clknet_leaf_82_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_69_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06930_ _02546_ _02564_ _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I spi_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06861_ _02330_ _02450_ _02496_ _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_08600_ ci_neuron.value_i\[22\] _03971_ _04078_ _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_06792_ _01892_ _02428_ _02429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_124_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05812_ _00739_ _01473_ _01474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09580_ net244 _04771_ _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05743_ _01359_ _01394_ _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08531_ ci_neuron.value_i\[12\] _04019_ _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05674_ _01223_ _01267_ _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08462_ ci_neuron.value_i\[2\] _03944_ net165 _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07413_ _02967_ _02968_ _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_64_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08393_ net529 net436 _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07344_ _02918_ _02920_ _02972_ _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_128_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout6_I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07275_ _01929_ _01937_ _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_115_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_135_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06226_ _01849_ _01859_ _01875_ _01876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04852__I _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09014_ _04361_ ci_neuron.stream_o\[8\] _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_135_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06157_ _01810_ _01811_ _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold131 ci_neuron.input_memory\[1\]\[3\] net555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold120 _04426_ net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold153 ci_neuron.output_val_internal\[27\] net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold142 ci_neuron.output_val_internal\[23\] net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_06088_ _01705_ _01718_ _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05108_ _00787_ _00770_ _00788_ _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold186 ci_neuron.output_val_internal\[26\] net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold175 ci_neuron.uut_simple_neuron.titan_id_6\[4\] net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold164 _00545_ net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold197 ci_neuron.input_memory\[1\]\[7\] net556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09916_ _00013_ net5 ci_neuron.address_i\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05039_ _00724_ _00725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09353__A2 _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09847_ _00426_ clknet_leaf_90_sys_clock_i ci_neuron.output_memory\[15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05914__A2 _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09778_ _00357_ clknet_leaf_139_sys_clock_i internal_ih.byte3\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_29_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08729_ _04187_ _04188_ _00587_ _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_96_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05602__A1 _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07355__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05390_ _01048_ _01051_ _01061_ _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__08607__A1 _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07060_ _02688_ _02692_ _02693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_3_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06011_ ci_neuron.uut_simple_neuron.x2\[27\] ci_neuron.uut_simple_neuron.x2\[28\]
+ _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05841__A1 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06397__A2 _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07594__A1 _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07962_ ci_neuron.uut_simple_neuron.titan_id_2\[22\] net458 _03533_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09701_ net3 clknet_leaf_103_sys_clock_i spi_interface_cvonk.MOSI_r\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold289_I ci_neuron.output_memory\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06913_ _02502_ _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07893_ ci_neuron.uut_simple_neuron.titan_id_2\[10\] net667 _03476_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06844_ _02057_ _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09632_ ci_neuron.stream_o\[18\] net261 _04811_ _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09563_ _04768_ _04769_ _04770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06775_ _02411_ _02356_ _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_104_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08514_ net124 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_104_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05726_ _01338_ _01340_ _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09494_ ci_neuron.output_memory\[18\] _04698_ _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_2_sys_clock_i_I clknet_4_1_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05657_ _01288_ _01294_ _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_77_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08445_ _03725_ _03945_ _03946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05588_ _01254_ _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08376_ _03880_ _03883_ _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07327_ _02954_ _02955_ _02956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04883__A2 _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07258_ _02886_ _02887_ _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07189_ _02819_ _02815_ _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06209_ ci_neuron.uut_simple_neuron.x3\[2\] _01859_ _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_103_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09865__CLK net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09574__A2 _04778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07888__A2 ci_neuron.uut_simple_neuron.titan_id_5\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09637__I0 ci_neuron.stream_o\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05588__I _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09262__A1 _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_23_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_90_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07328__A1 _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04890_ internal_ih.byte4\[2\] _00625_ _00628_ internal_ih.byte0\[2\] _00631_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_126_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06560_ _02200_ _02201_ _02202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_32_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_143_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06491_ _02099_ _02104_ _02133_ _02134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05511_ _01098_ _01150_ _01180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05442_ _01082_ _01112_ _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08230_ _03755_ _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_119_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05373_ _00939_ _01007_ _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08161_ net535 ci_neuron.uut_simple_neuron.titan_id_0\[27\] _03698_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_31_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07112_ _02380_ _02547_ _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08092_ net703 _00069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07043_ _02552_ _02624_ _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_2_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_41_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08994_ _04346_ _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07319__A1 _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07945_ _03517_ net484 _03519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_131_sys_clock_i clknet_4_2_0_sys_clock_i clknet_leaf_131_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07876_ net564 net304 _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09615_ ci_neuron.stream_o\[11\] net325 _04800_ _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06827_ _02401_ _02404_ _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_143_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06758_ _02395_ _02396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09546_ ci_neuron.output_memory\[26\] _04744_ _04755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05709_ _01145_ _01333_ _01372_ _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09477_ _04596_ _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06689_ _02289_ _02292_ _02327_ _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_109_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08428_ _00724_ _03924_ _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08359_ _03868_ _00183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05805__A1 _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10252_ _00150_ clknet_leaf_4_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[30\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10183_ _00081_ clknet_leaf_15_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07730__A1 ci_neuron.uut_simple_neuron.titan_id_4\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06297__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold708 _03415_ net741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold719 _00977_ net752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05991_ _01607_ _01630_ _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07730_ ci_neuron.uut_simple_neuron.titan_id_4\[15\] ci_neuron.uut_simple_neuron.titan_id_3\[15\]
+ _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_137_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04942_ _00662_ _00015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07661_ _03279_ _03281_ _03282_ _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_04873_ internal_ih.byte4\[5\] internal_ih.byte3\[5\] _00601_ _00619_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06612_ _02166_ _02251_ _02252_ _02253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07592_ _02933_ _03012_ _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09400_ _03740_ ci_neuron.input_memory\[1\]\[4\] _00768_ _01874_ _04622_ _04623_
+ _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_36_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06543_ _02094_ _02142_ _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_88_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09331_ _04566_ _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06474_ _02117_ _00230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09262_ _04166_ _04138_ _04127_ _04536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout22_I net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05425_ ci_neuron.uut_simple_neuron.x2\[15\] _01096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08213_ net749 _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09193_ _03967_ _04496_ _04497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_126_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05356_ _01027_ _01028_ _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08144_ _03680_ net643 _03683_ _03684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_43_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05287_ _00864_ _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08075_ _03606_ _03615_ _03626_ _03627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_70_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09428__I _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07026_ _02128_ _02603_ _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04860__I _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09529__A2 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold24 net597 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold46 net795 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08977_ net385 _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold35 spi_interface_cvonk.SS_r\[1\] net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07960__A1 _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold57 net810 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07928_ net660 _00135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold68 ci_neuron.uut_simple_neuron.titan_id_6\[25\] net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold79 _00525_ net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07859_ net731 net539 _03447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09529_ _04724_ _04740_ _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08512__I0 _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09465__A1 ci_neuron.output_memory\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10235_ _00131_ clknet_leaf_86_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10166_ _00092_ clknet_leaf_84_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10097_ _00163_ clknet_leaf_61_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_85_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_106_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_139_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04945__I _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06190_ _01820_ _01840_ _01841_ _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05210_ _00886_ _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05141_ _00743_ _00798_ _00820_ _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_13_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold527 _03633_ net560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold505 internal_ih.received_byte_count\[4\] net651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold516 internal_ih.spi_rx_byte_i\[0\] net549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_123_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold549 _03349_ net582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_05072_ _00755_ _00160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold538 _03513_ net571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_115_Left_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08900_ net270 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09880_ _00040_ net20 ci_neuron.value_i\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08831_ _04122_ net480 _04210_ _04253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_127_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05974_ _01601_ _01632_ _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08762_ _03955_ _04209_ _04213_ _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07713_ ci_neuron.uut_simple_neuron.titan_id_4\[12\] net677 _03327_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08498__A2 _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08693_ net238 _04137_ _04157_ _04155_ _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_04925_ _00639_ _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07644_ _03263_ _03266_ _03268_ _03269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_79_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_124_Left_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08528__S _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04856_ _00597_ _00602_ _00606_ internal_ih.byte7\[0\] _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_07575_ _02081_ _02480_ _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06526_ _02125_ _02128_ _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09314_ _04046_ net73 _04567_ _04569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06457_ _01963_ _01880_ _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09245_ _04526_ _00469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_145_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05408_ _01038_ _01062_ _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06388_ _02030_ _02016_ _02032_ _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09176_ _04484_ _00442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05339_ _00812_ _00847_ _00867_ _01011_ _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_08127_ _03670_ _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05236__A2 _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08058_ _03611_ net562 _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_56_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07009_ _02519_ _02518_ _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10020_ net77 clknet_leaf_19_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_1_0_sys_clock_i clknet_0_sys_clock_i clknet_4_1_0_sys_clock_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_85_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05475__A2 _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04986__A1 internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10218_ _00115_ clknet_leaf_31_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07924__A1 _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10149_ _00214_ clknet_leaf_38_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09516__I2 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05690_ _01353_ _01354_ _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_77_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08575__C _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07360_ _02986_ _02987_ _02910_ _02978_ _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_128_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06311_ _01957_ _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07291_ _02897_ _02908_ _02919_ _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_116_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09030_ _04377_ _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06242_ _01825_ _01852_ _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_143_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06173_ _01825_ _01822_ _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold302 _04294_ net335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05124_ _00786_ _00802_ _00803_ _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold313 _04329_ net346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold324 internal_ih.byte5\[6\] net357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold335 _04815_ net368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05055_ _00739_ _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold357 net830 net390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09932_ _00447_ clknet_leaf_76_sys_clock_i ci_neuron.uut_simple_neuron.x0\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold368 _04335_ net401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold346 ci_neuron.stream_o\[16\] net379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold379 _03315_ net412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08168__A1 _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09863_ _00442_ clknet_leaf_2_sys_clock_i ci_neuron.output_memory\[31\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08814_ _04085_ _01433_ _04239_ _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_51_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09794_ _00373_ clknet_leaf_137_sys_clock_i internal_ih.byte5\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08745_ net209 _04199_ internal_ih.received_byte_count\[5\] _04201_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05957_ _01614_ _01615_ _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05888_ _01548_ _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_107_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08676_ net125 _04137_ _04142_ _04143_ _04144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_04908_ _00642_ _00023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_138_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07627_ _03157_ _03193_ _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04839_ _00583_ internal_ih.received_byte_count\[2\] _00585_ _00590_ _00591_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07558_ _03182_ _03183_ _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06509_ _02130_ _02151_ _02152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07489_ _03109_ _03115_ _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08643__A2 _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09228_ _04059_ _03841_ _04514_ _04517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_51_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09159_ net102 _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08520__I _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10003_ net56 clknet_leaf_82_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05393__A1 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06645__A1 _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_93_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09673__D _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09526__I _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06860_ _02494_ _02495_ _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05811_ _01472_ _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06791_ _01983_ _02009_ _02428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_124_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05742_ _01405_ _00213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08530_ _04000_ _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_05673_ _01103_ _01332_ _01337_ _01338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_77_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08461_ _03735_ _03958_ _03959_ _03960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07412_ _03039_ _02998_ _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_135_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08392_ _03897_ _00187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07343_ _02962_ _02971_ _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_102_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07274_ _01920_ _02903_ _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold401_I internal_ih.byte7\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06225_ _01872_ _01874_ _01875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_14_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09013_ _04357_ _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_135_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold110 _00522_ net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_130_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06156_ _01615_ _01766_ _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold121 _00407_ net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold143 _00539_ net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold132 _03960_ net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06087_ _01741_ _01742_ _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05107_ _00773_ _00757_ _00768_ _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_hold770_I internal_ih.byte1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold176 net651 net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold154 _00543_ net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold165 net627 net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold198 net33 net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09915_ _00011_ net14 ci_neuron.address_i\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05038_ _00722_ _00723_ _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold187 _00542_ net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09846_ _00425_ clknet_leaf_88_sys_clock_i ci_neuron.output_memory\[14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07364__A2 _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08561__A1 _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06989_ ci_neuron.uut_simple_neuron.x3\[21\] _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05375__A1 _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09777_ _00356_ clknet_leaf_139_sys_clock_i internal_ih.byte3\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08728_ _04178_ net26 _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_1_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08313__A1 _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08659_ spi_interface_cvonk.state\[2\] spi_interface_cvonk.state\[1\] _04127_ _04128_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_96_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09041__A2 ci_neuron.stream_o\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05669__A2 ci_neuron.uut_simple_neuron.x2\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09655__I1 net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09668__D _00255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06010_ _01667_ _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07043__A1 _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_130_sys_clock_i clknet_4_2_0_sys_clock_i clknet_leaf_130_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07961_ net525 _00141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06912_ _02500_ _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09700_ net68 clknet_leaf_104_sys_clock_i spi_interface_cvonk.SS_r\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07892_ net669 _00128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06843_ _02477_ _02478_ _02479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09631_ net277 _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09591__I0 ci_neuron.stream_o\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06774_ _02411_ _02356_ _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09562_ _03904_ ci_neuron.input_memory\[1\]\[28\] _01792_ _03230_ _04760_ _04761_
+ _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA_hold449_I internal_ih.byte3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05725_ _01218_ _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05109__A1 _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08513_ _04004_ _00259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09343__I0 _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09493_ _04697_ _04707_ _04709_ _04710_ _00533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05656_ _00888_ _01174_ _01320_ _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_93_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08444_ _03942_ _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_137_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05587_ _01212_ _01253_ _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08375_ _03881_ _03882_ _03883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07326_ _02332_ _02882_ _02955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_92_sys_clock_i_I clknet_4_11_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07257_ _01908_ _02828_ _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07188_ _02282_ _02818_ _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06208_ ci_neuron.uut_simple_neuron.x3\[3\] ci_neuron.uut_simple_neuron.x3\[4\] _01859_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_115_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06139_ _01792_ _01793_ _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_112_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_6_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05596__A1 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08534__A1 _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05348__A1 _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09829_ _00408_ clknet_leaf_107_sys_clock_i internal_ih.spi_tx_byte_o\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09334__I0 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09262__A2 _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_56_sys_clock_i clknet_4_15_0_sys_clock_i clknet_leaf_56_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_90_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08773__A1 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09951__D _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09573__I0 _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09325__I0 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06490_ _02131_ _02132_ _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05510_ _00858_ _01178_ _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_136_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05441_ _01108_ _01111_ _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05511__A1 _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08160_ _03692_ _03695_ _03696_ _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09628__I1 ci_neuron.output_memory\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07111_ _02724_ _02742_ _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05372_ _01042_ _01019_ _01043_ _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08091_ _03639_ net702 _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07042_ _02672_ _02673_ _02674_ _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05814__A2 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09005__A2 _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07016__A1 _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__04873__I0 internal_ih.byte4\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08764__A1 _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08993_ net286 _04340_ _04346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_76_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07944_ ci_neuron.uut_simple_neuron.titan_id_2\[20\] net483 _03518_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07875_ _03453_ _03459_ _03460_ _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06826_ _02462_ _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_80_sys_clock_i_I clknet_4_14_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09614_ net356 _00561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09316__I0 _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04858__I _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06757_ _02135_ _02394_ _02395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09545_ _04743_ _04751_ _04753_ _04754_ _00541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06688_ _02282_ _02326_ _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05708_ _01191_ _01335_ _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_19_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09476_ _04673_ _04690_ _04694_ _04695_ _00531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05639_ _01240_ _01278_ _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05502__A1 _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08427_ _03925_ _03926_ _03927_ _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_47_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08358_ _03862_ _03864_ _03867_ _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_18_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07309_ _02937_ ci_neuron.uut_simple_neuron.x3\[25\] _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08289_ net621 _00174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10251_ _00148_ clknet_leaf_2_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05569__A1 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10182_ _00080_ clknet_leaf_15_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_141_Right_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold709 ci_neuron.uut_simple_neuron.titan_id_1\[25\] net742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_40_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_108_sys_clock_i_I clknet_4_9_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05990_ _01449_ _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04941_ internal_ih.byte6\[6\] _00658_ _00659_ internal_ih.byte2\[6\] _00662_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_88_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07660_ ci_neuron.uut_simple_neuron.titan_id_4\[3\] ci_neuron.uut_simple_neuron.titan_id_3\[3\]
+ _03282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_04872_ _00618_ _00029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07591_ _03148_ _03149_ _03212_ _03216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06611_ _02167_ _02207_ _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05732__A1 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06542_ _02045_ net274 _02183_ _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_88_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09330_ _04577_ _00503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09261_ _04534_ _04184_ _04124_ _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09474__A2 _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06473_ _02070_ _02116_ _02117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08212_ net174 _03740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05424_ _00860_ _01090_ _01094_ _01095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_90_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09192_ _04487_ _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout15_I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05355_ _00993_ _00994_ _01026_ _01028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08143_ net642 ci_neuron.uut_simple_neuron.titan_id_0\[23\] _03683_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_141_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08074_ _03614_ _03617_ _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08985__A1 _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07025_ _02606_ _02632_ _02657_ _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05286_ _00935_ _00946_ _00947_ _00949_ _00959_ _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_30_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_112_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold47 net804 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09444__I _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold25 net626 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_54_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08976_ net384 internal_ih.byte6\[5\] _04332_ _04336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold36 ci_neuron.uut_simple_neuron.x0\[0\] net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_145_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07927_ _03502_ _03503_ _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold58 net805 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold69 ci_neuron.uut_simple_neuron.titan_id_6\[23\] net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_97_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07858_ _03442_ _03445_ _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07789_ _03389_ _00112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06809_ _02383_ _02445_ _02446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_94_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09528_ _03864_ ci_neuron.input_memory\[1\]\[23\] _01433_ _02928_ _04738_ _04739_
+ _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__08512__I1 _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07476__A1 _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09459_ _04673_ _04676_ _04679_ _04681_ _00528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_136_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_27_sys_clock_i_I clknet_4_6_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07139__I _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10234_ _00130_ clknet_leaf_59_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10165_ _00091_ clknet_leaf_83_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10096_ _00162_ clknet_leaf_63_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09878__CLK net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_4_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09456__A2 _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05140_ _00735_ _00813_ _00816_ _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_52_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold517 ci_neuron.uut_simple_neuron.x2\[20\] net550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold506 ci_neuron.uut_simple_neuron.titan_id_5\[6\] net539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_122_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05071_ _00752_ _00754_ _00755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold528 ci_neuron.uut_simple_neuron.titan_id_1\[9\] net561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold539 _03514_ net572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08830_ _04252_ _00328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05973_ _01604_ _01631_ _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08761_ _00745_ _04211_ _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_127_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07712_ _03322_ _03324_ _03325_ _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_04924_ _00651_ _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08692_ _04141_ _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07643_ _03176_ _03179_ _03267_ _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04855_ _00605_ _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_140_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05705__B2 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07574_ _03198_ _03199_ _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09313_ _04568_ _00495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08608__I _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09447__A2 _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06525_ _02073_ _02159_ _02158_ _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_119_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07458__A1 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06456_ _01876_ _02100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09244_ _04094_ _03893_ _04525_ _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05407_ _00959_ _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_90_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09175_ net182 _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06387_ _02013_ _02031_ net54 _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08126_ net664 net778 _03670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05338_ _00983_ _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_4_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05269_ _00941_ _00943_ _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08057_ net561 ci_neuron.uut_simple_neuron.titan_id_0\[9\] _03612_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_56_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07008_ _02576_ _02588_ _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05944__A1 _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08959_ _04326_ _00383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_15_sys_clock_i_I clknet_4_1_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09438__A2 _04662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_80_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09461__I2 _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10217_ _00114_ clknet_leaf_40_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10148_ _00213_ clknet_leaf_38_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10079_ _00176_ clknet_leaf_118_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09516__I3 _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06360__A1 _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07290_ _02852_ _02896_ _02919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_128_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06310_ _01868_ _01934_ _01956_ _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06241_ _01889_ _01863_ _01885_ _01890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_142_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05787__I _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06172_ ci_neuron.uut_simple_neuron.x3\[0\] _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05123_ _00789_ _00799_ _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold314 ci_neuron.uut_simple_neuron.x0\[14\] net347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold325 _04328_ net358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold303 ci_neuron.stream_o\[9\] net336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05054_ _00738_ _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold369 ci_neuron.uut_simple_neuron.x0\[22\] net402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold336 net808 net369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold358 internal_ih.byte4\[2\] net391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold347 _04812_ net380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09931_ _00446_ clknet_leaf_77_sys_clock_i ci_neuron.uut_simple_neuron.x0\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold381_I ci_neuron.uut_simple_neuron.titan_id_5\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09862_ _00441_ clknet_leaf_2_sys_clock_i ci_neuron.output_memory\[30\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08813_ _04079_ _04211_ _04243_ _00320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_51_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _00372_ clknet_leaf_136_sys_clock_i internal_ih.byte5\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05956_ _01327_ _01478_ _01524_ _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_08744_ _04194_ _04200_ _00294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08539__S _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04907_ internal_ih.byte5\[0\] _00640_ _00641_ internal_ih.byte1\[0\] _00642_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05887_ _01511_ _01512_ _01546_ _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_107_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08675_ net549 _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07626_ _03249_ _03250_ _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04838_ _00586_ _00588_ _00589_ _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07557_ _02082_ _03113_ _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06508_ _02134_ _02150_ _02151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_75_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07488_ _03112_ _03114_ _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06439_ _02081_ _02082_ _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09227_ _04516_ _00461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09158_ _04475_ _00433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08109_ net589 _00072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09089_ ci_neuron.output_val_internal\[29\] ci_neuron.output_val_internal\[21\] ci_neuron.output_val_internal\[13\]
+ ci_neuron.output_val_internal\[5\] _04366_ _04367_ _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08651__I0 ci_neuron.uut_simple_neuron.x0\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08801__I _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10002_ net90 clknet_leaf_80_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_69_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_143_Left_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05810_ ci_neuron.uut_simple_neuron.x2\[24\] _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06790_ _02425_ _02426_ _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_124_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05741_ _01400_ _01404_ _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05672_ _01336_ _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08460_ _03942_ _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_07411_ _03028_ _03038_ _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08391_ _03890_ _03892_ _03896_ _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07342_ _02963_ _02970_ _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07273_ _01895_ _01899_ _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06224_ _01873_ _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09012_ internal_ih.data_pointer\[0\] _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_135_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06155_ _01613_ _01765_ _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold100 ci_neuron.uut_simple_neuron.titan_id_6\[15\] net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_130_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05106_ _00781_ _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold122 ci_neuron.uut_simple_neuron.titan_id_6\[16\] net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold133 ci_neuron.output_val_internal\[20\] net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold111 ci_neuron.output_val_internal\[16\] net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold144 ci_neuron.output_val_internal\[5\] net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06086_ _01412_ _01697_ _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold177 _04201_ net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold166 _00544_ net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold155 ci_neuron.output_val_internal\[21\] net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold188 internal_ih.received_byte_count\[0\] net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09914_ _00010_ net11 ci_neuron.address_i\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05037_ ci_neuron.address_i\[1\] ci_neuron.address_i\[0\] ci_neuron.address_i\[2\]
+ _00723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold199 ci_neuron.uut_simple_neuron.titan_id_6\[28\] net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09845_ _00424_ clknet_leaf_85_sys_clock_i ci_neuron.output_memory\[13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08936__I1 internal_ih.byte4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06988_ _02616_ _02556_ _02621_ _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_29_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09776_ _00355_ clknet_leaf_0_sys_clock_i internal_ih.byte3\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09452__I _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05939_ _01597_ _01598_ _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_68_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08727_ _04177_ _04186_ _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_29_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08313__A2 _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08658_ net404 _04127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07609_ _03168_ _03169_ _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_64_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08589_ _04011_ _04069_ _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04886__A1 internal_ih.byte4\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04886__B2 internal_ih.byte0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09577__A1 ci_neuron.output_memory\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_55_sys_clock_i clknet_4_15_0_sys_clock_i clknet_leaf_55_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_9_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09362__I _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06315__A1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08441__I _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07960_ _03530_ _03531_ _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_130_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06911_ _02505_ _02508_ _02545_ _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07891_ _03473_ _03474_ _03475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06842_ _02040_ _02437_ _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09272__I _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09630_ ci_neuron.stream_o\[17\] net276 _04811_ _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_136_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06773_ _02355_ _02411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09561_ _04700_ _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05724_ _01369_ _01387_ _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08512_ _04003_ _02089_ _03969_ _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09492_ net134 _04705_ _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05655_ _01083_ _01210_ _01176_ _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_77_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08443_ _03943_ _03944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_137_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05586_ _00860_ _01207_ _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08374_ _03869_ _03872_ _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07325_ _02341_ _02881_ _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07256_ _02273_ _02291_ _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06207_ _01821_ _01843_ _01839_ _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_60_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07187_ net318 _02817_ _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06580__B _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07034__A2 _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06138_ net746 _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06069_ _01594_ _01725_ _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05596__A2 _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09828_ net154 clknet_leaf_107_sys_clock_i internal_ih.spi_tx_byte_o\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09759_ _00338_ clknet_leaf_130_sys_clock_i internal_ih.byte1\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09098__I0 ci_neuron.output_val_internal\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08845__I0 internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05339__A2 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05440_ _01109_ _01110_ _01061_ _01059_ _01008_ _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
Xclkbuf_4_9_0_sys_clock_i clknet_0_sys_clock_i clknet_4_9_0_sys_clock_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09089__I0 ci_neuron.output_val_internal\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05371_ _01002_ _01011_ _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05511__A2 _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07110_ _02739_ _02741_ _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_119_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05275__A1 _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08090_ net701 ci_neuron.uut_simple_neuron.titan_id_0\[14\] _03640_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07041_ _02619_ _02627_ _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08992_ _04345_ _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold294_I ci_neuron.output_memory\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07943_ _03515_ _03516_ _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06527__A1 _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07874_ ci_neuron.uut_simple_neuron.titan_id_2\[7\] ci_neuron.uut_simple_neuron.titan_id_5\[7\]
+ ci_neuron.uut_simple_neuron.titan_id_2\[6\] net539 _03460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_06825_ _02418_ _02461_ _02462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09613_ net355 ci_neuron.output_memory\[10\] _04800_ _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06756_ _02096_ _02230_ _02394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_09544_ net225 _04749_ _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06687_ _02182_ _02287_ _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05707_ _01188_ _01370_ _01104_ _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_78_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09475_ net109 _04680_ _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05638_ _01300_ _01303_ _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_65_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08426_ _00709_ _03923_ _00728_ _00714_ _03927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_93_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05569_ _01169_ _01197_ _01237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08827__I0 _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08357_ _03865_ _03866_ _03867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07308_ ci_neuron.uut_simple_neuron.x3\[26\] _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08288_ _03803_ _03806_ _03807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07239_ _02868_ ci_neuron.uut_simple_neuron.x3\[24\] _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_132_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09252__I0 _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10250_ _00147_ clknet_leaf_3_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10181_ _00079_ clknet_leaf_17_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07191__A1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04940_ _00661_ _00014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__04959__I _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04871_ internal_ih.byte7\[4\] _00616_ _00617_ _00610_ _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07590_ _03215_ _00248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06610_ _02167_ _02207_ _02251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06541_ _02181_ _02182_ _02183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_87_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06472_ _02072_ _02115_ _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09260_ spi_interface_cvonk.SS_r\[2\] _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_16_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05423_ _01018_ _01093_ _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08211_ ci_neuron.uut_simple_neuron.x0\[4\] _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08682__A1 _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09191_ _03961_ _04494_ _04495_ _00446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05354_ _00993_ _00994_ _01026_ _01027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_83_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08142_ net644 _00079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05285_ _00879_ _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08073_ net674 _00095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07024_ _02608_ _02631_ _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06748__A1 _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09872__D _00063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08975_ net401 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_145_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07926_ ci_neuron.uut_simple_neuron.titan_id_2\[17\] ci_neuron.uut_simple_neuron.titan_id_5\[17\]
+ _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold26 ci_neuron.input_memory\[1\]\[8\] net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold37 spi_interface_cvonk.SCLK_r\[1\] net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold59 net803 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold48 ci_neuron.input_memory\[1\]\[23\] net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_98_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07857_ _03443_ _03444_ _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07788_ net446 net781 _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06808_ _02388_ _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_97_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06739_ _02332_ _02341_ _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09527_ _04668_ _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08673__A1 _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09458_ net127 _04680_ _04681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08409_ ci_neuron.uut_simple_neuron.x0\[28\] net417 _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09389_ net122 _04600_ _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06739__A1 _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08728__A2 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10233_ _00129_ clknet_leaf_88_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10164_ _00090_ clknet_leaf_83_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10095_ net97 clknet_leaf_61_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09370__I _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05190__A3 _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06978__A1 _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold507 _03450_ net540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold518 ci_neuron.uut_simple_neuron.x0\[31\] net551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_05070_ _00733_ net767 _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold529 _03612_ net562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05972_ _01607_ _01630_ _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08760_ _03947_ _04209_ _04212_ _00298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_29_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_127_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07155__A1 _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07711_ ci_neuron.uut_simple_neuron.titan_id_4\[11\] ci_neuron.uut_simple_neuron.titan_id_3\[11\]
+ _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08691_ _04134_ net118 _04156_ _00285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04923_ internal_ih.byte5\[7\] _00646_ _00647_ internal_ih.byte1\[7\] _00651_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07642_ _03162_ _03174_ _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04854_ _00604_ _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_140_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07573_ _03109_ _03115_ _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09312_ _04040_ net87 _04567_ _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06524_ _02119_ _02163_ _02165_ _02166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05469__A1 _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07458__A2 _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08825__S _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06455_ _02098_ _02088_ _02099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_118_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09243_ _04487_ _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_17_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06386_ _01947_ _01971_ _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05406_ _01076_ _01064_ _01077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09455__I0 _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09174_ _04483_ _00441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05337_ _01006_ _01008_ _01009_ _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08125_ ci_neuron.uut_simple_neuron.titan_id_1\[20\] net777 _03669_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_44_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05268_ _00909_ _00942_ _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08056_ _03609_ _03610_ _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07007_ _02637_ _02640_ _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05199_ _00876_ _00226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_47_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08430__I1 _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08958_ net430 net421 _04322_ _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07146__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07909_ _03485_ _03487_ _03488_ _03489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08889_ net489 net509 _04285_ _04287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09446__I0 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09461__I3 _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10216_ _00113_ clknet_leaf_40_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[26\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09365__I _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10147_ _00212_ clknet_leaf_43_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10078_ _00175_ clknet_leaf_71_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_122_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06240_ _01857_ _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_127_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09437__I0 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06171_ _01824_ _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_124_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07612__A2 _03233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05122_ _00789_ _00799_ _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold315 _03808_ net348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold304 _04802_ net337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold326 internal_ih.byte2\[5\] net359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05053_ ci_neuron.uut_simple_neuron.x2\[1\] _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05623__A1 _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold337 _04274_ net370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold359 _04313_ net392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold348 internal_ih.spi_rx_byte_i\[7\] net381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09930_ _00445_ clknet_leaf_77_sys_clock_i ci_neuron.uut_simple_neuron.x0\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09861_ _00440_ clknet_leaf_2_sys_clock_i ci_neuron.output_memory\[29\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08812_ _01381_ _04221_ _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09792_ _00371_ clknet_leaf_144_sys_clock_i internal_ih.byte5\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05955_ _01580_ _01613_ _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05308__I _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08743_ net209 _04199_ _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_84_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04906_ _00627_ _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05886_ _01511_ _01512_ _01546_ _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_89_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08674_ _04141_ _04142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07625_ _02121_ _03204_ _03250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04837_ internal_ih.expected_byte_count\[3\] _00584_ internal_ih.received_byte_count\[5\]
+ internal_ih.received_byte_count\[1\] _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07556_ _02489_ _02507_ _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_66_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06507_ _02147_ _02149_ _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_24_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07487_ _02082_ _03113_ _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07300__A1 _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09226_ _04052_ _03840_ _04514_ _04516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06438_ _02053_ _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07851__A2 ci_neuron.uut_simple_neuron.titan_id_5\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06369_ _02014_ _02012_ _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09157_ net257 _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_54_sys_clock_i clknet_4_15_0_sys_clock_i clknet_leaf_54_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_82_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08108_ net588 _03654_ _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09088_ _04417_ ci_neuron.stream_o\[5\] ci_neuron.stream_o\[21\] _04418_ _04430_
+ _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_141_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08039_ ci_neuron.uut_simple_neuron.titan_id_1\[6\] ci_neuron.uut_simple_neuron.titan_id_0\[6\]
+ _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_55_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10001_ net79 clknet_leaf_79_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_64_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_88_sys_clock_i_I clknet_4_11_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_136_Right_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05740_ _01313_ _01401_ _01403_ _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08439__I _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05671_ _01333_ _01335_ _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07410_ _03031_ _03037_ _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08390_ _03894_ _03895_ _03896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07341_ _02966_ _02969_ _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_9_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07272_ _02900_ _02901_ _02902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06223_ ci_neuron.uut_simple_neuron.x3\[4\] _01873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09011_ internal_ih.data_pointer\[1\] internal_ih.data_pointer\[0\] _04359_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_135_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06154_ _01756_ _01759_ _01808_ _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold101 ci_neuron.output_val_internal\[17\] net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05105_ _00779_ _00785_ _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold134 _00536_ net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold112 _00532_ net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold123 ci_neuron.output_val_internal\[13\] net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_06085_ _01557_ _01696_ _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold167 internal_ih.spi_tx_byte_o\[4\] net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold156 _00537_ net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold145 _00521_ net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold189 _00443_ net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold178 _00295_ net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09913_ _00009_ net7 ci_neuron.address_i\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05036_ ci_neuron.address_i\[22\] ci_neuron.address_i\[23\] _00716_ _00721_ _00722_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09844_ _00423_ clknet_leaf_85_sys_clock_i ci_neuron.output_memory\[12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_119_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06987_ _02551_ _02620_ _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09775_ _00354_ clknet_leaf_0_sys_clock_i internal_ih.byte3\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05938_ _01547_ _01552_ _01548_ _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08726_ _04178_ _04183_ _04185_ _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_29_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05869_ _01529_ _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08657_ spi_interface_cvonk.SCLK_r\[2\] _04125_ _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07608_ _03231_ _03232_ _03233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08588_ _03996_ _04067_ _04068_ _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_48_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07539_ _03163_ _03164_ _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09209_ _04506_ _00453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_122_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07856__C ci_neuron.uut_simple_neuron.titan_id_5\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_92_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold690 _03510_ net723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_76_sys_clock_i_I clknet_4_10_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06315__A2 _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09265__A1 _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_145_sys_clock_i_I clknet_4_0_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06910_ _02497_ _02504_ _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07890_ ci_neuron.uut_simple_neuron.titan_id_2\[10\] net667 _03474_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09553__I _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06841_ _02041_ _02436_ _02477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07751__A1 _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06772_ _02406_ _02409_ _02410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09560_ net198 _04766_ _04767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05723_ _01374_ _01378_ _01386_ _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_78_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08511_ _03996_ _03998_ _03999_ _04002_ _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_09491_ _04701_ _04708_ _04709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07503__A1 _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08442_ _03942_ _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05654_ _01318_ _01296_ _01297_ _01284_ _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_93_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05585_ _01179_ _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08373_ _03863_ net388 _03881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07324_ _02951_ _02952_ _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07255_ _02855_ _02884_ _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_61_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06206_ _01856_ _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09875__D _00035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07186_ _02441_ _02740_ _02816_ _02817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_112_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06137_ _01668_ _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06068_ _01691_ _01724_ _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_6_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05019_ net170 _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09827_ net217 clknet_leaf_106_sys_clock_i internal_ih.spi_tx_byte_o\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08790__I0 _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09758_ _00337_ clknet_leaf_130_sys_clock_i internal_ih.byte0\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08709_ _04167_ net184 _04130_ _00290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09689_ _00276_ clknet_leaf_26_sys_clock_i ci_neuron.uut_simple_neuron.x3\[26\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05339__A3 _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09238__A1 _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_133_sys_clock_i_I clknet_4_2_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05370_ _01039_ _01040_ _01041_ _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_16_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07040_ _02629_ _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_11_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08452__I _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09410__A1 ci_neuron.output_memory\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08991_ _04155_ net530 _04339_ _04345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_76_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07942_ _03512_ _03513_ _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07873_ _03457_ _03458_ _03459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06824_ _02422_ _02460_ _02461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09612_ net337 _00560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09543_ _04746_ _04752_ _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_143_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06755_ _02382_ _02392_ _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_78_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06686_ _01928_ _02324_ _02325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_93_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05706_ _01191_ _01335_ _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_19_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09474_ _04677_ _04693_ _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05637_ _01078_ _01301_ _01302_ _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08425_ _00708_ _00709_ ci_neuron.stream_enabled _03923_ _03926_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_2
X_08356_ _03856_ _03859_ _03866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05568_ _00959_ _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07307_ _02928_ _02869_ _02935_ _02936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05499_ _01134_ _01155_ _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08287_ _03804_ _03805_ _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_61_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07238_ ci_neuron.uut_simple_neuron.x3\[25\] _02868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07169_ ci_neuron.uut_simple_neuron.x3\[23\] ci_neuron.uut_simple_neuron.x3\[24\]
+ _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_76_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09252__I1 _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10180_ _00078_ clknet_leaf_17_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07963__A1 _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09368__I _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_121_sys_clock_i_I clknet_4_3_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04870_ internal_ih.byte4\[4\] internal_ih.byte3\[4\] _00608_ _00617_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08648__S _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06540_ _02144_ _02182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_88_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06471_ _02114_ _02112_ _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05422_ _00982_ _01092_ _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08210_ _03738_ _00194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08682__A2 _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09190_ _03724_ _04491_ _04495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05353_ _00996_ _01025_ _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_83_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08141_ _03680_ net643 _03682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05284_ _00953_ _00956_ _00951_ _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08072_ _03623_ net673 _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07023_ _01857_ _02655_ _02656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_58_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08974_ net400 internal_ih.byte6\[4\] _04332_ _04335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_145_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06430__I _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold27 net628 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07925_ _03500_ _03501_ _03502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold38 net753 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_145_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold49 ci_neuron.output_memory\[2\] net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_07856_ ci_neuron.uut_simple_neuron.titan_id_2\[5\] ci_neuron.uut_simple_neuron.titan_id_5\[5\]
+ ci_neuron.uut_simple_neuron.titan_id_2\[4\] ci_neuron.uut_simple_neuron.titan_id_5\[4\]
+ _03444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07787_ net780 ci_neuron.uut_simple_neuron.titan_id_3\[25\] _03388_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06807_ _02280_ _02391_ _02443_ _02444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_04999_ internal_ih.byte2\[7\] _00691_ _00695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06738_ _01958_ _02375_ _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09526_ _04666_ _04738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__04931__A1 internal_ih.byte6\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09457_ _04610_ _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06669_ _02301_ _02307_ _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08408_ _03903_ _03905_ _03911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_81_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09388_ _04598_ _04617_ _04619_ _04620_ _00518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_47_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08339_ _03850_ _03851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_40_sys_clock_i_I clknet_4_5_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06987__A2 _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06739__A2 _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10232_ _00128_ clknet_leaf_87_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10163_ _00089_ clknet_leaf_83_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09528__I2 _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10094_ _00192_ clknet_leaf_5_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08267__I _03788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06978__A2 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold508 _03452_ net541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold519 internal_ih.byte0\[4\] net552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_122_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05971_ _01567_ _01629_ _01630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07710_ ci_neuron.uut_simple_neuron.titan_id_4\[11\] ci_neuron.uut_simple_neuron.titan_id_3\[11\]
+ _03324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_53_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04922_ _00650_ _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08690_ _04155_ _04149_ _04156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07641_ _03264_ _03189_ _03265_ _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04853_ _00594_ _00603_ _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_140_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07572_ _03112_ _03114_ _03198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_109_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06523_ _02120_ _02162_ _02165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09311_ _04566_ _04567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__04913__B2 internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06454_ net230 _02097_ _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09242_ _04524_ _00468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08905__I _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06385_ _02018_ _02019_ _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05405_ _01075_ _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09173_ net179 _04483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05336_ _00852_ _00972_ _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08124_ net663 ci_neuron.uut_simple_neuron.titan_id_0\[19\] _03657_ _03665_ _03667_
+ _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xclkbuf_leaf_53_sys_clock_i clknet_4_15_0_sys_clock_i clknet_leaf_53_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_102_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05267_ _00914_ _00942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08055_ _03606_ _03607_ _03610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07006_ _02638_ _02573_ _02639_ _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_141_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05198_ _00851_ _00875_ _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07394__A2 _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08957_ net424 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07908_ net473 ci_neuron.uut_simple_neuron.titan_id_5\[13\] _03488_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09471__I _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08888_ _04286_ _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07839_ net608 ci_neuron.uut_simple_neuron.titan_id_5\[3\] _03429_ _03430_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_84_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09509_ _04700_ _04724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_137_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10215_ _00112_ clknet_leaf_40_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_120_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07166__I ci_neuron.uut_simple_neuron.x3\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10146_ _00211_ clknet_leaf_43_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05396__A1 _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10077_ _00174_ clknet_leaf_71_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_46_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06170_ _01823_ _01824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05121_ _00801_ _00223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold316 ci_neuron.uut_simple_neuron.x3\[31\] net349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold305 ci_neuron.input_memory\[1\]\[30\] net338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05052_ _00736_ _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold349 _04266_ net382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold327 _04295_ net360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold338 ci_neuron.stream_o\[13\] net371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09860_ _00439_ clknet_leaf_1_sys_clock_i ci_neuron.output_memory\[28\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05387__A1 _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08811_ _04242_ _00319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09791_ _00370_ clknet_leaf_144_sys_clock_i internal_ih.byte5\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05954_ _01326_ _01612_ _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08742_ _04193_ net272 _04199_ _00293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_108_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08673_ _04138_ _04140_ _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_04905_ _00639_ _00640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07624_ _02131_ _02103_ _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05885_ _01076_ _01545_ _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_95_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_04836_ internal_ih.expected_byte_count\[0\] _00587_ _00588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07555_ _03159_ _03180_ _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07486_ _02489_ _02507_ _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_119_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06506_ _01925_ _02148_ _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06437_ _02047_ _02081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07300__A2 _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09225_ _04515_ _00460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06368_ _01947_ _01971_ _02013_ _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09156_ _04474_ _00432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_142_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06299_ _01867_ _01936_ _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05319_ _00992_ _00203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08107_ _03653_ _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09087_ _04405_ _04429_ _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08038_ net690 _00090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_2_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10000_ net86 clknet_leaf_79_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05378__A1 _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09989_ _00504_ clknet_leaf_11_sys_clock_i ci_neuron.input_memory\[1\]\[24\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06802__A1 _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09376__I _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10129_ _00161_ clknet_leaf_61_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_124_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06869__A1 _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05670_ _01226_ _01290_ _01334_ _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09107__I0 ci_neuron.output_val_internal\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07340_ _02967_ _02968_ _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_128_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07271_ _02824_ _02830_ _02901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09010_ _04357_ _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06222_ _01838_ _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06153_ _01714_ _01760_ _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05104_ _00780_ _00754_ _00782_ _00784_ _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
Xhold113 ci_neuron.uut_simple_neuron.titan_id_6\[17\] net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold102 _00533_ net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold135 ci_neuron.output_val_internal\[7\] net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold124 _00529_ net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_06084_ _01738_ _01739_ _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold168 _04160_ net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold157 net687 net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold146 ci_neuron.uut_simple_neuron.titan_id_6\[30\] net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05319__I _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold179 ci_neuron.uut_simple_neuron.x0\[6\] net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_10_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05035_ _00717_ _00718_ _00719_ _00720_ _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_09912_ _00008_ net7 ci_neuron.address_i\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09843_ _00422_ clknet_leaf_89_sys_clock_i ci_neuron.output_memory\[11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06986_ _02555_ _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09774_ _00353_ clknet_leaf_0_sys_clock_i internal_ih.byte2\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05937_ _01593_ _01596_ _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_68_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08725_ _04184_ _04140_ _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05868_ _01479_ _01525_ _01529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08656_ net70 _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_139_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07607_ _03229_ _03230_ ci_neuron.uut_simple_neuron.x3\[29\] _03232_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08587_ ci_neuron.value_i\[20\] _04055_ _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07538_ _02870_ _03091_ _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05799_ _01377_ _01371_ _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07469_ _03094_ _03095_ _03096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09208_ _04003_ _03772_ _04488_ _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_79_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09139_ net151 _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08785__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold680 ci_neuron.uut_simple_neuron.titan_id_4\[2\] net713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_9_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold691 ci_neuron.uut_simple_neuron.titan_id_1\[10\] net724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09585__I0 _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05771__A1 _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09265__A2 _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08776__A1 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10192__D _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06840_ _01847_ _02428_ _02475_ _02476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_65_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06771_ _02309_ _02407_ _02408_ _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05762__A1 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05722_ _01384_ _01385_ _01386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09490_ _03824_ ci_neuron.input_memory\[1\]\[17\] _01184_ _02445_ _04691_ _04692_
+ _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08510_ ci_neuron.value_i\[9\] _04001_ _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05653_ _01286_ _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08441_ _03925_ _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05584_ _01215_ _01249_ _01250_ _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_63_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08372_ net389 _03879_ _03880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07323_ _01948_ _02892_ _02952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_83_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07254_ _02883_ _02879_ _02884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06205_ _01852_ _01854_ _01855_ _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_104_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04876__I0 internal_ih.byte4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07185_ _02442_ _02615_ _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06136_ _01789_ _01767_ _01790_ _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06067_ _01650_ _01723_ _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_41_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05018_ _00705_ _00057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08519__A1 ci_neuron.value_i\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_92_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09826_ _00405_ clknet_leaf_106_sys_clock_i internal_ih.spi_tx_byte_o\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06969_ _02173_ _02148_ _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08790__I1 _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09757_ _00336_ clknet_leaf_130_sys_clock_i internal_ih.byte0\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08708_ net183 _04168_ _04131_ _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09688_ _00275_ clknet_leaf_26_sys_clock_i ci_neuron.uut_simple_neuron.x3\[25\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05505__A1 _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08639_ _04110_ _03230_ _04111_ _04112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout30 net31 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07430__A1 _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09573__I3 ci_neuron.uut_simple_neuron.x3\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05744__A1 _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05339__A4 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08990_ _04170_ _04340_ _04344_ _00396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09564__I _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07972__A2 net624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07941_ ci_neuron.uut_simple_neuron.titan_id_2\[19\] ci_neuron.uut_simple_neuron.titan_id_5\[19\]
+ _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07872_ _03447_ _03451_ _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06823_ _02424_ _02459_ _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09611_ net336 ci_neuron.output_memory\[9\] _04800_ _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06754_ _02391_ _02280_ _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09542_ _03893_ ci_neuron.input_memory\[1\]\[25\] _01573_ _02934_ _04738_ _04739_
+ _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_143_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05705_ _01341_ _01346_ _01367_ _01368_ _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA_hold447_I ci_neuron.uut_simple_neuron.x2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06685_ _01935_ _02323_ _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09473_ _03825_ ci_neuron.input_memory\[1\]\[15\] _01098_ _02387_ _04691_ _04692_
+ _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_19_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05636_ _01251_ _01275_ _01302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08424_ _00724_ _03924_ _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_46_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05567_ _01067_ _01234_ _01235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10097__D _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08355_ _03850_ net291 _03865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07306_ _02863_ _02934_ _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_34_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05498_ _01134_ _01155_ _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08286_ _03783_ _03796_ _03794_ _03805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_33_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07237_ _02731_ _02864_ _02866_ _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_33_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07168_ _02734_ _02735_ _02798_ _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_76_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06119_ _01771_ _01774_ _01775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07099_ _02730_ _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09809_ _00388_ clknet_leaf_136_sys_clock_i internal_ih.byte7\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08818__I _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_145_sys_clock_i clknet_4_0_0_sys_clock_i clknet_leaf_145_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_122_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06390__A1 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06470_ _02113_ _02063_ _02114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_16_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05421_ _00964_ _01055_ _01091_ _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_16_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08140_ net642 ci_neuron.uut_simple_neuron.titan_id_0\[23\] _03681_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05352_ _00905_ _01024_ _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05283_ _00957_ _00202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08071_ net672 ci_neuron.uut_simple_neuron.titan_id_0\[11\] _03624_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07022_ _02653_ _02654_ _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold397_I internal_ih.byte6\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08973_ net398 _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_145_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07924_ _03497_ _03498_ _03501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold28 net556 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_145_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold39 net714 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07855_ ci_neuron.uut_simple_neuron.titan_id_2\[5\] ci_neuron.uut_simple_neuron.titan_id_5\[5\]
+ _03443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07786_ net445 ci_neuron.uut_simple_neuron.titan_id_3\[24\] _03376_ _03384_ _03386_
+ _03387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_06806_ _02441_ _02442_ _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05184__A2 _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08638__I _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04998_ _00694_ _00047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06737_ _02374_ _01968_ _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09525_ ci_neuron.output_memory\[23\] _04722_ _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06668_ _02250_ _02253_ _02302_ _02304_ _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_78_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09456_ _04677_ _04678_ _04679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05619_ _01262_ _01271_ _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08407_ _03905_ net647 _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06599_ _02219_ _02221_ _02239_ _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09387_ ci_neuron.output_val_internal\[2\] _04611_ _04620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08338_ net429 _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07633__A1 _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09473__I2 _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08269_ _03782_ _03784_ _03778_ _03779_ _03777_ _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_6_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10231_ _00158_ clknet_leaf_85_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10162_ _00088_ clknet_leaf_83_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10093_ _00191_ clknet_leaf_5_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[30\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09528__I3 _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold509 ci_neuron.uut_simple_neuron.x0\[16\] net542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05970_ _01628_ _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_53_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04921_ internal_ih.byte5\[6\] _00646_ _00647_ internal_ih.byte1\[6\] _00650_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_127_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07640_ _03184_ _03191_ _03265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04852_ _00599_ _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_140_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07571_ _03195_ _03196_ _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_109_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06522_ _02164_ _00231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09310_ _04542_ _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06453_ _02093_ _02096_ _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_75_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09241_ _04089_ _03877_ _04519_ _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06706__I _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06384_ _01945_ _02021_ _02028_ _02015_ _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_05404_ _01067_ _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout13_I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09172_ _04482_ _00440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05335_ _00964_ _01007_ _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08123_ _03660_ _03666_ _03667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08054_ ci_neuron.uut_simple_neuron.titan_id_1\[8\] ci_neuron.uut_simple_neuron.titan_id_0\[8\]
+ _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07005_ _02569_ _02572_ _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_114_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05266_ _00938_ _00940_ _00941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05197_ _00854_ _00874_ _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA_hold779_I ci_neuron.uut_simple_neuron.titan_id_5\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08956_ internal_ih.byte6\[4\] net423 _04322_ _04325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07907_ ci_neuron.uut_simple_neuron.titan_id_2\[13\] ci_neuron.uut_simple_neuron.titan_id_5\[13\]
+ _03487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08887_ net466 net502 _04285_ _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06354__A1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07838_ _03425_ _03427_ _03428_ _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_116_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07769_ net640 ci_neuron.uut_simple_neuron.titan_id_3\[22\] _03372_ _03373_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_84_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09508_ ci_neuron.output_memory\[20\] _04722_ _04723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09439_ net113 _04655_ _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10214_ _00111_ clknet_leaf_41_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_95_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10145_ _00210_ clknet_leaf_43_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10076_ _00173_ clknet_leaf_72_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_122_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08893__I0 internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09437__I2 _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05120_ _00778_ _00800_ _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08645__I0 _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold306 internal_ih.byte6\[1\] net339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold317 ci_neuron.normalised_stream_write_address\[0\] net350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05051_ _00735_ _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold339 _04807_ net372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold328 ci_neuron.output_memory\[31\] net361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_41_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07357__I _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08810_ _04074_ _01368_ _04239_ _04242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08573__A2 _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09790_ _00369_ clknet_leaf_144_sys_clock_i internal_ih.byte4\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05953_ ci_neuron.uut_simple_neuron.x2\[23\] _01379_ _01524_ _01612_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08741_ net271 _04197_ _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05884_ _01515_ _01544_ _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_04904_ _00604_ _00639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08672_ net300 _04139_ _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07623_ _03246_ _03247_ _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04898__A1 internal_ih.byte4\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_04835_ net221 _00587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07554_ _03176_ _03179_ _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_119_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04898__B2 internal_ih.byte0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07485_ _03110_ _03111_ _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06505_ _01905_ _02000_ _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06436_ _01833_ _02079_ _02080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_90_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09224_ _04046_ _03822_ _04514_ _04515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06367_ _01951_ _01970_ _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_90_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09155_ net251 _04474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06298_ _01944_ _01940_ _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05318_ _00958_ _00991_ _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_82_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08106_ ci_neuron.uut_simple_neuron.titan_id_1\[17\] ci_neuron.uut_simple_neuron.titan_id_0\[17\]
+ _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09086_ _04419_ ci_neuron.stream_o\[13\] _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05249_ _00885_ _00923_ _00924_ _00901_ _00855_ _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_08037_ net689 _03594_ _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_130_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09988_ _00503_ clknet_leaf_30_sys_clock_i ci_neuron.input_memory\[1\]\[23\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08939_ _04315_ _00374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_103_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08875__I0 internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06802__A2 _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_112_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10128_ _00160_ clknet_leaf_62_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_124_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10059_ net199 clknet_leaf_123_sys_clock_i ci_neuron.output_val_internal\[28\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_121_Left_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06869__A2 _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05541__A2 _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08866__I0 internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07270_ _02827_ _02829_ _02900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06221_ _01870_ _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_135_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_130_Left_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06152_ _01648_ _01806_ _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08471__I _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06083_ _01604_ _01723_ _01739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05103_ _00783_ _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold125 internal_ih.expected_byte_count\[2\] net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold114 internal_ih.spi_tx_byte_o\[5\] net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold103 ci_neuron.output_val_internal\[19\] net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_112_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09911_ _00007_ net7 ci_neuron.address_i\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05034_ ci_neuron.address_i\[9\] ci_neuron.address_i\[8\] ci_neuron.address_i\[7\]
+ ci_neuron.address_i\[6\] _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold158 _04395_ net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold147 ci_neuron.output_val_internal\[0\] net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold136 _00523_ net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_112_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold169 _00287_ net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold477_I internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09842_ _00421_ clknet_leaf_88_sys_clock_i ci_neuron.output_memory\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09773_ _00352_ clknet_leaf_0_sys_clock_i internal_ih.byte2\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06985_ _02442_ _02558_ _02618_ _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08724_ spi_interface_cvonk.SCLK_r\[2\] _04125_ _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05936_ _01594_ _01545_ _01595_ _01596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_68_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05867_ _01477_ _01479_ _01480_ _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08655_ net68 _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07606_ _03229_ _03230_ _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08586_ _03848_ _04066_ _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_clkbuf_leaf_129_sys_clock_i_I clknet_4_2_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05532__A2 _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07537_ _03087_ _03089_ _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05798_ _01458_ _01459_ _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07468_ _02682_ _02930_ _03095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08482__A1 _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07399_ _03004_ _03021_ _03026_ _03027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06419_ _02029_ _02033_ _02063_ _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__08609__I0 _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09207_ _03994_ _04503_ _04505_ _00452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09138_ _04465_ _00423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09477__I _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09069_ internal_ih.spi_tx_byte_o\[3\] _04379_ _04414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06260__A3 _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold670 _03641_ net703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold681 ci_neuron.input_memory\[1\]\[25\] net775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_9_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold692 _03619_ net725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__05220__A1 _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_101_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_48_sys_clock_i_I clknet_4_6_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06770_ _02351_ _02353_ _02408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05721_ _00740_ _01343_ _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05652_ _01075_ _01299_ _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08440_ _03940_ _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_81_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05583_ _01217_ _01231_ _01250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_63_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08371_ _03878_ _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07322_ _02323_ _02344_ _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold225_I ci_neuron.output_val_internal\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07253_ _02332_ _02882_ _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_128_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07184_ _02796_ _02811_ _02814_ _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_121_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06204_ _01825_ _01845_ _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_54_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04876__I1 internal_ih.byte3\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06135_ _01753_ _01761_ _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06066_ _01694_ _01722_ _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_117_sys_clock_i_I clknet_4_9_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05017_ internal_ih.byte3\[7\] _00701_ _00705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08519__A2 _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09825_ _00404_ clknet_leaf_106_sys_clock_i internal_ih.spi_tx_byte_o\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06968_ _02600_ _02601_ _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09756_ _00335_ clknet_leaf_105_sys_clock_i internal_ih.byte0\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09687_ _00274_ clknet_leaf_27_sys_clock_i ci_neuron.uut_simple_neuron.x3\[24\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05919_ ci_neuron.uut_simple_neuron.x2\[26\] _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08707_ _04166_ _04141_ _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06899_ _02532_ _02533_ _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08638_ _03939_ _04111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08569_ _03968_ _04053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_65_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09952__CLK clknet_4_4_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout31 internal_ih.got_all_data net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout20 net21 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_144_sys_clock_i clknet_4_0_0_sys_clock_i clknet_leaf_144_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_33_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09089__I3 ci_neuron.output_val_internal\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08446__A1 ci_neuron.value_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_36_sys_clock_i_I clknet_4_5_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_51_sys_clock_i clknet_4_13_0_sys_clock_i clknet_leaf_51_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_31_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09246__I0 _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05680__A1 _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05594__B _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05432__A1 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07940_ net572 _00137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07871_ _03455_ _03456_ _03445_ _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06822_ _02431_ _02458_ _02459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09610_ net352 _00559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06753_ _02386_ _02390_ _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09541_ ci_neuron.output_memory\[25\] _04744_ _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05704_ _01344_ _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06684_ _02044_ _02290_ _02322_ _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09472_ _04668_ _04692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_19_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05635_ _01251_ _01275_ _01301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_19_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08423_ _00714_ _03923_ _00710_ _03924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05566_ _01206_ _01233_ _01234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08354_ _03863_ _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_105_sys_clock_i_I clknet_4_8_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07305_ _02868_ _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05497_ _01164_ _01165_ _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08285_ _03794_ ci_neuron.uut_simple_neuron.x0\[13\] _03790_ _03791_ _03789_ _03804_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_6_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07236_ _02797_ _02865_ _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_15_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07167_ _02730_ _02797_ _02798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_76_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06118_ _01772_ _01773_ _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07098_ ci_neuron.uut_simple_neuron.x3\[22\] _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06049_ ci_neuron.uut_simple_neuron.x2\[27\] _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07176__A1 _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09808_ _00387_ clknet_leaf_0_sys_clock_i internal_ih.byte7\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09739_ _00318_ clknet_leaf_30_sys_clock_i ci_neuron.uut_simple_neuron.x2\[20\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08676__B2 _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09228__I0 _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08600__A1 ci_neuron.value_i\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_24_sys_clock_i_I clknet_4_6_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05420_ _00969_ ci_neuron.uut_simple_neuron.x2\[13\] ci_neuron.uut_simple_neuron.x2\[14\]
+ _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_127_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05351_ _00999_ _01023_ _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_44_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05282_ _00954_ _00956_ _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_70_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08070_ _03621_ _03622_ _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09219__I0 _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07021_ _02599_ _02605_ _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08972_ net397 internal_ih.byte6\[3\] _04332_ _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold292_I ci_neuron.output_memory\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07923_ net645 net659 _03500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold29 net666 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_145_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold557_I ci_neuron.uut_simple_neuron.titan_id_5\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07854_ _03434_ _03435_ _03440_ _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06805_ _02387_ _02389_ _02442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_39_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07785_ _03385_ _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_04997_ internal_ih.byte2\[6\] _00691_ _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06736_ _02085_ _02343_ _02373_ _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_94_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09524_ _04721_ _04733_ _04735_ _04736_ _00538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06667_ _02306_ _00234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09455_ _03795_ ci_neuron.input_memory\[1\]\[12\] _00971_ _02226_ _04667_ _04669_
+ _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
Xclkbuf_leaf_19_sys_clock_i clknet_4_6_0_sys_clock_i clknet_leaf_19_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05618_ _01260_ _01284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08406_ _03909_ _00189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06598_ _02235_ _02238_ _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09386_ _04603_ _04618_ _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05549_ _01183_ _01194_ _01216_ _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08337_ _03848_ _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09473__I3 _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08268_ net366 net386 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__08425__A4 _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07219_ _02792_ _02832_ _02849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10230_ _00157_ clknet_leaf_86_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08199_ net528 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09485__I _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07397__A1 _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10161_ _00077_ clknet_leaf_91_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10092_ _00189_ clknet_leaf_6_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08821__A1 _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_12_sys_clock_i_I clknet_4_4_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09377__A2 _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04920_ _00649_ _00005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_127_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07560__A1 _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04851_ internal_ih.byte4\[0\] internal_ih.byte3\[0\] _00601_ _00602_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_140_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06259__I _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07570_ _00162_ _03129_ _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_7_sys_clock_i_I clknet_4_4_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06521_ _02119_ _02163_ _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_109_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09240_ _04523_ _00467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06452_ _02001_ _02095_ _02096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_91_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06383_ _02018_ _02019_ _02028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05403_ _01032_ _01063_ _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09171_ net237 _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05334_ _00970_ _01006_ _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08812__A1 _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09455__I3 _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08122_ ci_neuron.uut_simple_neuron.titan_id_1\[19\] ci_neuron.uut_simple_neuron.titan_id_0\[19\]
+ _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08053_ net656 _00092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07004_ _02515_ _02517_ _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_141_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05265_ _00939_ _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_131_Right_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05196_ _00855_ _00873_ _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08955_ _04324_ _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07906_ net474 _00131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08886_ _04269_ _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_98_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_16_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07837_ ci_neuron.uut_simple_neuron.titan_id_2\[2\] ci_neuron.uut_simple_neuron.titan_id_5\[2\]
+ _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07768_ _03368_ net576 _03371_ _03372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06719_ _02308_ _02357_ _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_84_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09507_ _04674_ _04722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07699_ net411 ci_neuron.uut_simple_neuron.titan_id_3\[9\] _03312_ _03313_ _03315_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_94_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09438_ _04652_ _04662_ _04663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_81_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09369_ _03930_ _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_136_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08803__A1 _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09446__I3 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07606__A2 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_25_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05093__A2 _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10213_ _00110_ clknet_leaf_42_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_120_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10144_ _00209_ clknet_leaf_42_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10075_ _00172_ clknet_leaf_72_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_34_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07845__A2 net590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09437__I3 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold307 _04331_ net340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06820__A3 _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05050_ _00734_ _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold329 ci_neuron.output_memory\[0\] net362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold318 ci_neuron.stream_o\[8\] net351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05952_ _00748_ _01582_ _01581_ _01610_ _01529_ _01611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_08740_ net271 _04197_ _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05883_ _01518_ _01520_ _01543_ _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_84_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08671_ net249 spi_interface_cvonk.state\[0\] _04139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_04903_ _00638_ _00022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09522__A2 _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09373__I2 _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07622_ _00163_ _03206_ _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04834_ internal_ih.received_byte_count\[4\] internal_ih.received_byte_count\[7\]
+ internal_ih.received_byte_count\[6\] _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_36_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07553_ _02550_ _03178_ _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09286__A1 _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07484_ _02444_ _03025_ _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06504_ _02138_ _02146_ _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_66_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06435_ _01868_ _01954_ _02078_ _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_107_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09223_ _04499_ _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_106_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09154_ _04473_ _00431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06366_ _01987_ _01993_ _02011_ _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08105_ _03648_ _03649_ _03651_ _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_16_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06297_ _01909_ _01911_ _01944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05317_ _00960_ _00990_ _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09085_ _04415_ net153 _04428_ _00407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05248_ _00889_ _00899_ _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08036_ ci_neuron.uut_simple_neuron.titan_id_1\[6\] ci_neuron.uut_simple_neuron.titan_id_0\[6\]
+ _03594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09210__A1 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05179_ _00835_ _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09987_ _00502_ clknet_leaf_72_sys_clock_i ci_neuron.input_memory\[1\]\[22\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08938_ net423 net428 _04312_ _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_4_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08869_ net502 net504 _04275_ _04276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09277__A1 _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05838__A1 _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10127_ _00159_ clknet_leaf_62_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_124_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10058_ net187 clknet_leaf_121_sys_clock_i ci_neuron.output_val_internal\[27\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07515__A1 _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09268__A1 _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05829__A1 _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06220_ _01867_ _01861_ _01869_ _01870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08491__A2 _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06151_ _01785_ _01788_ _01805_ _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_81_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06272__I _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06082_ _01694_ _01722_ _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05102_ _00734_ _00770_ _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold126 _00513_ net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold115 _04162_ net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold104 _00535_ net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold137 ci_neuron.uut_simple_neuron.x0\[1\] net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09910_ _00006_ net8 ci_neuron.address_i\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05033_ ci_neuron.address_i\[5\] ci_neuron.address_i\[4\] ci_neuron.address_i\[3\]
+ _00719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xhold148 _00516_ net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold159 ci_neuron.output_val_internal\[4\] net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09841_ _00420_ clknet_leaf_85_sys_clock_i ci_neuron.output_memory\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_119_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06984_ _02615_ _02617_ _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09772_ _00351_ clknet_leaf_1_sys_clock_i internal_ih.byte2\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05935_ _01515_ _01544_ _01595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08723_ _04179_ _04182_ _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_68_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05866_ _01526_ _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08654_ _04123_ _00281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05797_ _01437_ _01439_ _01459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07605_ net756 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08585_ _03838_ _04049_ _04066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_119_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07536_ _03160_ _03161_ _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07467_ _02727_ _02867_ _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09206_ _03770_ _04500_ _04505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_143_sys_clock_i clknet_4_0_0_sys_clock_i clknet_leaf_143_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_17_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07398_ _02444_ _03025_ _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06418_ _02062_ _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_20_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06349_ _01966_ _01995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09137_ net129 _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09431__A1 ci_neuron.output_memory\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06245__A1 _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09068_ net215 _04381_ _04412_ _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08019_ ci_neuron.uut_simple_neuron.titan_id_1\[2\] net287 _03580_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold660 ci_neuron.uut_simple_neuron.titan_id_4\[16\] net693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold671 ci_neuron.uut_simple_neuron.titan_id_4\[29\] net704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_120_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_9_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold682 _03279_ net715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold693 _03620_ net726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09881__CLK net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08793__I0 _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05220__A2 _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07741__I net582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05261__I _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_50_sys_clock_i clknet_4_13_0_sys_clock_i clknet_leaf_50_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_101_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05720_ _01329_ _01380_ _01383_ _01384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_78_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05651_ _01283_ _01298_ _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_4_12_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08370_ _03877_ _03875_ _03878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07321_ _02924_ _02949_ _02950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_129_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05582_ _01217_ _01231_ _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_63_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08839__I1 _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08464__A2 _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_69_sys_clock_i clknet_4_12_0_sys_clock_i clknet_leaf_69_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_144_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07252_ _02341_ _02881_ _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06203_ _01853_ _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07183_ _02494_ _02813_ _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_60_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07098__I ci_neuron.uut_simple_neuron.x3\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06134_ _01762_ _01789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06065_ _01699_ _01721_ _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_6_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05016_ _00704_ _00056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09824_ _00403_ clknet_leaf_110_sys_clock_i internal_ih.spi_tx_byte_o\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_4_6_0_sys_clock_i clknet_0_sys_clock_i clknet_4_6_0_sys_clock_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06967_ _02131_ _02543_ _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09755_ _00334_ clknet_leaf_132_sys_clock_i internal_ih.byte0\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06898_ _02047_ _02490_ _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09686_ _00273_ clknet_leaf_27_sys_clock_i ci_neuron.uut_simple_neuron.x3\[23\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05918_ _01472_ _01577_ _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08706_ internal_ih.spi_rx_byte_i\[7\] _04166_ _04142_ _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_139_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05849_ _01510_ _00215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08637_ _04107_ _04108_ _04109_ _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_139_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08568_ _04048_ _04050_ _04051_ _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_49_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout10 net15 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout21 net22 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07519_ _03143_ _03144_ _03145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08499_ _03769_ _03987_ _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xfanout32 net69 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08455__A2 _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold490 _03301_ net523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08766__I0 _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08391__A1 _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08694__A2 _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09246__I1 _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05432__A2 _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07870_ _03435_ _03440_ _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06821_ _02434_ _02457_ _02458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06752_ _02387_ _02389_ _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09540_ _04743_ _04745_ _04748_ _04750_ _00540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05703_ _00750_ _01329_ _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09471_ _04666_ _04691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06683_ _02045_ _02181_ _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_18_sys_clock_i clknet_4_3_0_sys_clock_i clknet_leaf_18_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08422_ ci_neuron.instruction_i\[2\] _03922_ _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_19_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05634_ _01067_ _01299_ _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05115__B _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05565_ _01215_ _01232_ _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08353_ net399 _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07304_ _02734_ _02735_ _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06448__A1 _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08284_ net620 net347 _03803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_46_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05496_ _01075_ _01157_ _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07235_ ci_neuron.uut_simple_neuron.x3\[24\] _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07166_ ci_neuron.uut_simple_neuron.x3\[23\] _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_76_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07097_ _02548_ _02683_ _02728_ _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06117_ _01699_ _01721_ _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06048_ _01663_ _01703_ _01704_ _01621_ _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_30_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07176__A2 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09807_ _00386_ clknet_leaf_140_sys_clock_i internal_ih.byte7\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07999_ net498 _03542_ _03559_ _03564_ _03565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_97_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09738_ _00317_ clknet_leaf_29_sys_clock_i ci_neuron.uut_simple_neuron.x2\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09669_ _00256_ clknet_4_13_0_sys_clock_i ci_neuron.uut_simple_neuron.x3\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_145_Right_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08987__I0 _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08600__A2 _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_129_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06678__A1 _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_16_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05350_ _01001_ _01004_ _01022_ _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_83_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05281_ _00927_ _00926_ _00928_ _00955_ _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_70_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07020_ _02602_ _02604_ _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08971_ net435 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_145_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07922_ _03499_ _00134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07158__A2 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07853_ net593 _00154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06804_ _02386_ _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_127_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07784_ ci_neuron.uut_simple_neuron.titan_id_4\[24\] ci_neuron.uut_simple_neuron.titan_id_3\[24\]
+ ci_neuron.uut_simple_neuron.titan_id_4\[23\] ci_neuron.uut_simple_neuron.titan_id_3\[23\]
+ _03385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_78_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_04996_ _00693_ _00046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06735_ _02086_ _02222_ _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09523_ net171 _04727_ _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06666_ _02303_ _02305_ _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_79_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09454_ _04602_ _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07330__A2 _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05617_ _01257_ _01274_ _01282_ _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09385_ _03724_ ci_neuron.input_memory\[1\]\[2\] _00774_ _01849_ _04605_ _04607_
+ _04618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08405_ _03904_ _03905_ _03908_ _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_19_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06597_ _02237_ _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08336_ ci_neuron.uut_simple_neuron.x0\[20\] _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05548_ _00751_ _01152_ _01193_ _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_34_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05479_ ci_neuron.uut_simple_neuron.x2\[16\] _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08267_ _03788_ _00171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07218_ _02792_ _02832_ _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_132_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06841__A1 _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_89_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08198_ _03728_ _00190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07149_ _02710_ _02711_ _02715_ _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_120_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07286__I _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08594__A1 _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10160_ _00066_ clknet_leaf_91_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10091_ _00188_ clknet_leaf_7_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_98_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04907__A1 internal_ih.byte5\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08821__A2 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10289_ _00582_ clknet_leaf_128_sys_clock_i ci_neuron.stream_o\[31\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04850_ _00600_ _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_140_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06520_ _02120_ _02162_ _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_109_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08755__I _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06451_ _02090_ _02094_ _02095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05402_ _01073_ _00205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05323__A1 _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06382_ _01981_ _02023_ _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_97_sys_clock_i_I clknet_4_10_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09170_ _04481_ _00439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05333_ _01005_ _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08121_ _03658_ _03663_ _03665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05264_ ci_neuron.uut_simple_neuron.x2\[9\] ci_neuron.uut_simple_neuron.x2\[10\]
+ ci_neuron.uut_simple_neuron.x2\[11\] _00939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_08052_ _03606_ net655 _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07003_ _02634_ _02636_ _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_114_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05195_ _00856_ _00872_ _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08954_ net444 net439 _04322_ _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07905_ net473 ci_neuron.uut_simple_neuron.titan_id_5\[13\] _03485_ _03486_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08885_ _04284_ _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09540__A3 _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07836_ ci_neuron.uut_simple_neuron.titan_id_2\[2\] ci_neuron.uut_simple_neuron.titan_id_5\[2\]
+ _03427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07767_ net575 ci_neuron.uut_simple_neuron.titan_id_3\[21\] _03371_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_04979_ _00683_ _00038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06718_ _02356_ _02355_ _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_84_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09506_ _04696_ _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07698_ net599 _00125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09701__D net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06649_ _02288_ _02282_ _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_109_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09437_ _04005_ net76 _00911_ _02091_ _04644_ _04645_ _04662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_13_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09368_ _04602_ _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09299_ net76 _04556_ _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08319_ net407 _03830_ _03831_ _03834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_145_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08803__A2 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10212_ _00109_ clknet_leaf_42_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_95_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10143_ _00208_ clknet_leaf_42_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10074_ _00171_ clknet_leaf_81_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06805__A1 _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08524__B _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold308 ci_neuron.stream_o\[12\] net341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold319 _04801_ net352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_55_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05951_ _01584_ _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_84_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_85_sys_clock_i_I clknet_4_14_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05882_ _01538_ _01542_ _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09373__I3 _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08670_ spi_interface_cvonk.SCLK_r\[2\] _04125_ _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_04902_ internal_ih.byte4\[7\] _00633_ _00634_ internal_ih.byte0\[7\] _00638_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07621_ _03203_ _03205_ _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04833_ _00583_ internal_ih.received_byte_count\[2\] internal_ih.expected_byte_count\[3\]
+ _00584_ _00585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07552_ _02559_ _03177_ _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06503_ _02045_ _02145_ _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_66_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07483_ _02451_ _03024_ _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_66_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06434_ _02055_ _02056_ _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09222_ _04513_ _00459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_57_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_142_sys_clock_i clknet_4_0_0_sys_clock_i clknet_leaf_142_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_17_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06365_ _02006_ _02010_ _02011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_56_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09153_ net243 _04473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05316_ _00879_ _00989_ _00990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08104_ ci_neuron.uut_simple_neuron.titan_id_1\[16\] ci_neuron.uut_simple_neuron.titan_id_0\[16\]
+ _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_114_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06296_ _01912_ _01914_ _01941_ _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09084_ internal_ih.spi_tx_byte_o\[4\] _04427_ _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05247_ _00889_ _00899_ _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08035_ _03590_ _03592_ _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05178_ _00820_ _00853_ _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09210__A2 _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09986_ _00501_ clknet_leaf_30_sys_clock_i ci_neuron.input_memory\[1\]\[21\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08937_ net440 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08868_ _04269_ _04275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07819_ net740 ci_neuron.uut_simple_neuron.titan_id_3\[30\] _03414_ _03415_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_4_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08799_ _04052_ net754 _04231_ _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09521__I0 _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06263__A2 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05259__I _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10126_ net231 clknet_leaf_62_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10057_ net220 clknet_leaf_128_sys_clock_i ci_neuron.output_val_internal\[26\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06818__I _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_68_sys_clock_i clknet_4_12_0_sys_clock_i clknet_leaf_68_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08779__A1 _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06150_ _01791_ _01804_ _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_73_sys_clock_i_I clknet_4_9_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06081_ _01736_ _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05101_ _00781_ _00761_ _00782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold116 _00288_ net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold105 ci_neuron.interrupt_enabled net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05032_ ci_neuron.address_i\[17\] ci_neuron.address_i\[16\] ci_neuron.address_i\[15\]
+ ci_neuron.address_i\[14\] _00718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold149 ci_neuron.uut_simple_neuron.titan_id_6\[31\] net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold127 ci_neuron.uut_simple_neuron.titan_id_6\[6\] net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold138 ci_neuron.output_val_internal\[22\] net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_42_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold198_I net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09840_ _00419_ clknet_leaf_88_sys_clock_i ci_neuron.output_memory\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06983_ _02616_ _02556_ _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09771_ _00350_ clknet_leaf_139_sys_clock_i internal_ih.byte2\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05934_ _01236_ _01594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08722_ _04173_ _04174_ _04181_ _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_68_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05865_ _01374_ _01461_ _01525_ _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08653_ _04122_ net349 _04111_ _04123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_135_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05796_ _01426_ _01457_ _01458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08584_ _04065_ _00269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07604_ net727 _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_53_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07535_ _03093_ _03097_ _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07466_ _03082_ _03092_ _03093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06417_ _01985_ _02036_ _02061_ _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_119_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09205_ _03990_ _04503_ _04504_ _00451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_142_sys_clock_i_I clknet_4_0_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04879__I0 internal_ih.byte4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07397_ _02451_ _03024_ _03025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_106_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06348_ _01963_ _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09136_ _04464_ _00422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06279_ _01925_ _01926_ _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_103_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09067_ _04382_ _04408_ _04410_ _04411_ _04412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_32_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08018_ net106 _00127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold672 _03411_ net705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold661 _03344_ net694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_92_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold650 ci_neuron.input_memory\[1\]\[21\] net761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_9_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold683 _03280_ net716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold694 _03084_ net727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09969_ _00484_ clknet_leaf_81_sys_clock_i ci_neuron.input_memory\[1\]\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05028__B _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06373__I _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07984__A2 net695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09186__A1 _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10109_ _00233_ clknet_leaf_53_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_61_sys_clock_i_I clknet_4_14_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05650_ _01315_ _00211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_17_sys_clock_i clknet_4_1_0_sys_clock_i clknet_leaf_17_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05581_ _01075_ _01234_ _01247_ _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07320_ _02945_ _02948_ _02949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_63_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08763__I _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07251_ _02494_ _02813_ _02880_ _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06202_ _01844_ _01853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07182_ _02449_ _02812_ _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06133_ _01786_ _01787_ _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08472__I0 _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07975__A2 ci_neuron.uut_simple_neuron.titan_id_5\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06064_ _01702_ _01720_ _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09177__B2 _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05015_ internal_ih.byte3\[6\] _00701_ _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_74_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09823_ _00402_ clknet_leaf_100_sys_clock_i internal_ih.instruction_received vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_130_sys_clock_i_I clknet_4_2_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06966_ _02132_ _02542_ _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09754_ _00333_ clknet_leaf_131_sys_clock_i internal_ih.byte0\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06897_ _02082_ _02489_ _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09685_ _00272_ clknet_leaf_24_sys_clock_i ci_neuron.uut_simple_neuron.x3\[22\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_05917_ ci_neuron.uut_simple_neuron.x2\[25\] ci_neuron.uut_simple_neuron.x2\[26\]
+ _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XPHY_EDGE_ROW_61_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08705_ _04147_ _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05848_ _01495_ _01509_ _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_96_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08636_ ci_neuron.value_i\[28\] _04001_ _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05779_ _01415_ _01441_ _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08567_ ci_neuron.value_i\[17\] _04032_ _04051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout11 net14 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout22 net23 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09101__A1 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07518_ _03066_ _03141_ _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08498_ _03986_ _03990_ _03991_ _00257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout33 ci_neuron.uut_simple_neuron.x2\[0\] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_134_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07449_ _03004_ _03021_ _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_33_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_70_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07415__A1 _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09119_ net247 _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05977__A1 _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold480 ci_neuron.uut_simple_neuron.titan_id_2\[30\] net513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_102_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08766__I1 _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold491 ci_neuron.uut_simple_neuron.titan_id_2\[22\] net524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08391__A2 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_109_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07957__A2 net414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_118_Left_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06820_ _02438_ _02440_ _02456_ _02457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__08758__I _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06751_ ci_neuron.uut_simple_neuron.x3\[16\] _02388_ _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_06682_ _02275_ _02294_ _02320_ _02321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05702_ _01362_ _01364_ _01365_ _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_78_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09470_ ci_neuron.output_memory\[15\] _04675_ _04690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08421_ _00711_ _00712_ _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05633_ _01283_ _01298_ _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09589__I _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_127_Left_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05564_ _01217_ _01231_ _01232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08352_ _03861_ _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_hold328_I ci_neuron.output_memory\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout29_I net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07303_ _02727_ net499 _02931_ _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__06448__A2 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05495_ _01126_ _01156_ _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08283_ _03802_ _00173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07234_ _02797_ _02863_ _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_143_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09398__A1 ci_neuron.output_memory\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07165_ _02739_ _02741_ _02795_ _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_76_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07096_ _02725_ _02727_ _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06116_ _01702_ _01720_ _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_136_Left_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06047_ _01668_ _01622_ _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09806_ _00385_ clknet_leaf_142_sys_clock_i internal_ih.byte6\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09570__A1 ci_neuron.output_val_internal\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07998_ net784 net618 _03558_ _03561_ _03563_ _03564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06949_ _02410_ _02357_ _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09737_ _00316_ clknet_leaf_26_sys_clock_i ci_neuron.uut_simple_neuron.x2\[18\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09668_ _00255_ clknet_leaf_65_sys_clock_i ci_neuron.uut_simple_neuron.x3\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_145_Left_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08619_ _04094_ _02934_ _04086_ _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09599_ _04789_ _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_77_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07747__I net712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09400__I2 _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05280_ _00922_ _00925_ _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06850__A2 _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08978__I1 internal_ih.byte6\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08970_ net434 internal_ih.byte6\[2\] _04332_ _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07921_ _03497_ net646 _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_71_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07852_ net592 _03440_ _03441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_hold180_I ci_neuron.output_val_internal\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold278_I ci_neuron.output_memory\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06803_ _02393_ _02396_ _02439_ _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xinput1 spi_clock_i net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07783_ _03377_ _03382_ _03384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_04995_ internal_ih.byte2\[5\] _00691_ _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09522_ _04724_ _04734_ _04735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06734_ _02325_ _02370_ _02371_ _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_hold445_I internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06665_ _02250_ _02253_ _02304_ _02305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09453_ ci_neuron.output_memory\[12\] _04675_ _04676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_143_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05616_ _01259_ _01273_ _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08404_ _03906_ _03907_ _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09384_ net82 _04600_ _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06596_ _01994_ _02236_ _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08335_ _03847_ _00180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05547_ _01105_ _01209_ _01182_ _01214_ _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_74_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05478_ _01097_ _01147_ _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_85_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08266_ _03782_ _03785_ net579 _03788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07217_ _02787_ _02788_ _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06841__A2 _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08197_ _03724_ _03727_ _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07148_ _02761_ _02763_ _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07079_ _02661_ _02667_ _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10090_ _00187_ clknet_leaf_9_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10288_ _00581_ clknet_leaf_128_sys_clock_i ci_neuron.stream_o\[30\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09534__A1 ci_neuron.output_memory\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06450_ ci_neuron.uut_simple_neuron.x3\[11\] _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05401_ _01071_ _01072_ _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_75_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_141_sys_clock_i clknet_4_0_0_sys_clock_i clknet_leaf_141_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08972__S _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06381_ _01981_ _02023_ _02025_ _02026_ _00228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_28_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05332_ ci_neuron.uut_simple_neuron.x2\[13\] _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08120_ net671 _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05263_ _00937_ _00916_ _00938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08051_ net654 ci_neuron.uut_simple_neuron.titan_id_0\[8\] _03607_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07002_ _02526_ _02568_ _02635_ _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_4_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05194_ _00841_ _00853_ _00871_ _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_40_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08953_ net450 _00380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07904_ _03481_ net377 _03484_ _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06339__A1 _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08884_ net359 net475 _04280_ _04284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05011__A1 internal_ih.byte3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07835_ net662 _00149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07766_ net577 _00108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04978_ internal_ih.byte1\[6\] _00680_ _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06717_ _02257_ _02299_ _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_84_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09505_ _04697_ _04715_ _04719_ _04720_ _00535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_07697_ _03312_ _03313_ _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09436_ ci_neuron.output_memory\[10\] _04650_ _04661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06648_ _02144_ _02287_ _02288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_109_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06579_ _02184_ _02190_ _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08639__I0 _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09367_ _00728_ _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09298_ _04559_ _00489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08318_ _03830_ _03831_ net407 _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_34_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08249_ _03756_ _03769_ _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10211_ _00108_ clknet_leaf_42_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_95_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10142_ _00207_ clknet_leaf_41_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10073_ _00170_ clknet_leaf_81_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_126_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05002__A1 internal_ih.byte3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_67_sys_clock_i clknet_4_12_0_sys_clock_i clknet_leaf_67_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_128_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold309 _04806_ net342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_33_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05950_ _01526_ _01586_ _01608_ _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05881_ _01252_ _01254_ _01541_ _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_04901_ _00637_ _00021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07620_ _03243_ _03244_ _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04832_ internal_ih.received_byte_count\[3\] _00584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07551_ _02725_ _03096_ _03095_ _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06502_ _02141_ _02144_ _02145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_88_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08869__I0 net502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07482_ _03107_ _03108_ _03109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06433_ _02039_ _02060_ _02076_ _02077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_91_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09221_ _04040_ _03825_ _04509_ _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06364_ _02009_ _02010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout11_I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09152_ _04472_ _00430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05315_ _00946_ _00988_ _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08103_ _03650_ _00071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06295_ _01942_ _00168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09083_ _04377_ _04427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05246_ _00905_ _00921_ _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08034_ _03588_ _03591_ _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05177_ _00735_ _00838_ _00833_ _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_12_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09985_ _00500_ clknet_leaf_26_sys_clock_i ci_neuron.input_memory\[1\]\[20\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08936_ net439 internal_ih.byte4\[3\] _04312_ _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08867_ net370 _00343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07818_ _03410_ _03412_ _03413_ _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_4_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06732__A1 _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08798_ _04234_ _00314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_109_sys_clock_i clknet_4_8_0_sys_clock_i clknet_leaf_109_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07749_ _03348_ _03353_ _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07288__A2 _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09521__I1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09419_ _04630_ _04646_ _04647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10125_ _00249_ clknet_leaf_35_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10056_ net226 clknet_leaf_122_sys_clock_i ci_neuron.output_val_internal\[25\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08712__A2 _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_16_sys_clock_i clknet_4_1_0_sys_clock_i clknet_leaf_16_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_106_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08476__A1 ci_neuron.value_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06080_ _01734_ _01735_ _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05100_ net33 _00781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xhold117 ci_neuron.uut_simple_neuron.titan_id_6\[10\] net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold106 ci_neuron.stream_o\[31\] net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_123_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold128 internal_ih.spi_tx_byte_o\[1\] net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05031_ ci_neuron.address_i\[13\] ci_neuron.address_i\[12\] ci_neuron.address_i\[11\]
+ ci_neuron.address_i\[10\] _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold139 _00538_ net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06982_ _02498_ _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09770_ _00349_ clknet_4_2_0_sys_clock_i internal_ih.byte2\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05933_ _01449_ _01592_ _01593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08721_ internal_ih.instruction_received internal_ih.spi_rx_byte_i\[3\] _04180_ _04181_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_68_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08652_ ci_neuron.value_i\[31\] _04121_ _04026_ _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07603_ _03226_ _03227_ _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05864_ _01327_ _01524_ _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_77_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05795_ _01432_ _01436_ _01457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_95_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08583_ _04064_ _02552_ _04053_ _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07534_ _03082_ _03092_ _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07465_ _02870_ _03091_ _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06416_ _02039_ _02060_ _02061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09204_ _03756_ _04500_ _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04879__I1 internal_ih.byte3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07396_ _02615_ _03022_ _03023_ _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_20_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06347_ _01989_ _01990_ _01992_ _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_115_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09135_ net205 _04464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06278_ _01905_ _01926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_79_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09066_ _04182_ _04411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05229_ _00787_ _00836_ _00904_ _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08017_ ci_neuron.uut_simple_neuron.titan_id_2\[0\] net105 _03579_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_92_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold662 ci_neuron.uut_simple_neuron.titan_id_5\[26\] net695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold640 _03624_ net673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold651 ci_neuron.uut_simple_neuron.titan_id_1\[26\] net684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold684 ci_neuron.uut_simple_neuron.titan_id_4\[23\] net717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_130_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold673 ci_neuron.uut_simple_neuron.titan_id_4\[11\] net706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__05205__A1 _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold695 ci_neuron.uut_simple_neuron.titan_id_5\[11\] net728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09195__A2 _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09968_ _00483_ clknet_4_12_0_sys_clock_i ci_neuron.input_memory\[1\]\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09578__S0 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08919_ internal_ih.byte4\[4\] net419 _04301_ _04304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09899_ _00018_ net9 ci_neuron.address_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09498__A3 _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05444__A1 _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07197__A1 _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09186__A2 _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10108_ _00232_ clknet_leaf_53_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10039_ net108 clknet_leaf_77_sys_clock_i ci_neuron.output_val_internal\[8\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05580_ _01206_ _01233_ _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_81_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08449__A1 _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07250_ _02495_ _02812_ _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08980__S _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06201_ _01842_ _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07181_ _02622_ _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07424__A2 _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06132_ _01450_ _01777_ _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05435__A1 _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08472__I1 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06063_ _01661_ _01719_ _01720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05014_ _00703_ _00054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_74_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09822_ _00401_ clknet_leaf_133_sys_clock_i internal_ih.current_instruction\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09753_ net228 clknet_leaf_132_sys_clock_i internal_ih.byte0\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06965_ _02597_ _02598_ _02599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08704_ _04133_ net131 _04165_ _00289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06896_ _02529_ _02530_ _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05916_ _00937_ _01575_ _01569_ _01576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09684_ _00271_ clknet_leaf_27_sys_clock_i ci_neuron.uut_simple_neuron.x3\[21\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08688__B2 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05847_ _01500_ _01502_ _01508_ _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08635_ _03904_ _04106_ _03959_ _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_138_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06163__A2 _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08566_ _03971_ _04049_ _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07517_ _03068_ _03140_ _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05778_ _01418_ _01440_ _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xfanout12 net14 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08497_ net824 _03980_ _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout23 net24 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07448_ _03028_ _03038_ _03074_ _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07379_ _03005_ _03006_ _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09118_ _04455_ _00413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09049_ net161 _04379_ _04396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold470 internal_ih.byte2\[0\] net503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold481 _03574_ net514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold492 _03532_ net525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_99_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05665__A1 _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06750_ ci_neuron.uut_simple_neuron.x3\[17\] _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06681_ _02278_ _02293_ _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05701_ _01331_ _01363_ _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07342__A1 _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05632_ _01284_ _01297_ _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08420_ _03921_ _00192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05563_ _01221_ _01230_ _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08351_ net402 _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05494_ _01163_ _00207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07302_ _02930_ _02870_ _02931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08282_ _03798_ _03801_ _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08842__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07233_ ci_neuron.uut_simple_neuron.x3\[24\] _02863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05656__A1 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07164_ _02729_ _02738_ _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_76_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07095_ _02726_ _02681_ _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06115_ _01698_ _01746_ _01770_ _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_30_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06046_ _01672_ _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__04919__B1 _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ _00384_ clknet_leaf_142_sys_clock_i internal_ih.byte6\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07997_ _03562_ _03563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06948_ _02578_ _02579_ _02580_ _02582_ _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_09736_ _00315_ clknet_leaf_24_sys_clock_i ci_neuron.uut_simple_neuron.x2\[17\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09667_ _00254_ clknet_leaf_65_sys_clock_i ci_neuron.uut_simple_neuron.x3\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06879_ _02472_ _02514_ _02515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_87_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08618_ _04091_ _04093_ _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_38_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09720__D _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07884__A2 ci_neuron.uut_simple_neuron.titan_id_5\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09598_ _04794_ _00554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08549_ _04035_ _00264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08617__C _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07636__A2 _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08859__I _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_5_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09400__I3 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05283__I _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_140_sys_clock_i clknet_4_0_0_sys_clock_i clknet_leaf_140_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07920_ net645 ci_neuron.uut_simple_neuron.titan_id_5\[16\] _03498_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07851_ ci_neuron.uut_simple_neuron.titan_id_2\[5\] ci_neuron.uut_simple_neuron.titan_id_5\[5\]
+ _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06802_ _02382_ _02392_ _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06366__A2 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07782_ net612 _00111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput2 spi_cs_i net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06733_ _02328_ _02346_ _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09521_ _03862_ net67 _01381_ _02805_ _04716_ _04717_ _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_04994_ _00692_ _00045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06664_ _02209_ _02249_ _02304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_94_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09452_ _04674_ _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05615_ _01281_ _00210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06595_ _01995_ _02093_ _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_08403_ _03898_ _03901_ _03907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09383_ _04598_ _04613_ _04615_ _04616_ _00517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_145_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05546_ _01212_ _01213_ _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08334_ _03844_ _03846_ _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05477_ _01146_ _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08265_ _03777_ _03780_ _03786_ _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07216_ _02835_ _02838_ _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08196_ _03725_ _03726_ _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07147_ _02774_ _02776_ _02777_ _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_104_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06054__A1 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07078_ _02664_ _02666_ _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06029_ _01686_ _00219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_89_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09543__A2 _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09719_ _00298_ clknet_leaf_67_sys_clock_i ci_neuron.uut_simple_neuron.x2\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_66_sys_clock_i clknet_4_13_0_sys_clock_i clknet_leaf_66_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10287_ _00580_ clknet_leaf_128_sys_clock_i ci_neuron.stream_o\[29\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09385__I2 _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07442__B _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07848__A2 net590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05400_ _01029_ _01027_ _01070_ _01072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_84_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06380_ _02024_ _02023_ _02026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05331_ _00743_ _01002_ _00974_ _01003_ _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_56_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09470__A1 ci_neuron.output_memory\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05262_ _00936_ _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05087__A2 _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08050_ _03602_ _03603_ _03604_ _03605_ _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_40_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07001_ _02528_ _02567_ _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05193_ _00862_ _00870_ _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08952_ internal_ih.byte6\[2\] net449 _04322_ _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07903_ ci_neuron.uut_simple_neuron.titan_id_2\[12\] net376 _03484_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08883_ _04283_ _00350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07834_ net661 ci_neuron.uut_simple_neuron.titan_id_5\[2\] _03425_ _03426_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_07765_ _03368_ net576 _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09289__A1 _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04977_ _00682_ _00037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_108_sys_clock_i clknet_4_9_0_sys_clock_i clknet_leaf_108_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06716_ _02309_ _02354_ _02355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07696_ net411 net598 _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_84_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09504_ net136 _04705_ _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06647_ _02285_ _02286_ _02287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_94_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08887__I1 net502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09435_ _04649_ _04657_ _04659_ _04660_ _00525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_93_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06578_ _01870_ _02218_ _02219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_118_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_69_sys_clock_i_I clknet_4_12_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08639__I1 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09366_ ci_neuron.output_memory\[0\] _04600_ _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_145_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05529_ _01169_ _01197_ _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09297_ _04003_ net58 _04543_ _04559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08317_ net406 ci_neuron.uut_simple_neuron.x0\[18\] _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08248_ _03771_ _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10210_ _00106_ clknet_leaf_44_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08179_ ci_neuron.uut_simple_neuron.titan_id_1\[29\] ci_neuron.uut_simple_neuron.titan_id_0\[29\]
+ _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_95_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10141_ _00206_ clknet_leaf_54_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10072_ _00199_ clknet_leaf_81_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_126_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_15_sys_clock_i clknet_4_1_0_sys_clock_i clknet_leaf_15_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_69_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_138_sys_clock_i_I clknet_4_2_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08878__I1 net481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07518__A1 _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04900_ internal_ih.byte4\[6\] _00633_ _00634_ internal_ih.byte0\[6\] _00637_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05880_ _01429_ _01539_ _01540_ _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_84_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_04831_ net158 _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07550_ _03175_ _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06501_ _02090_ _02143_ _02144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_07481_ _02041_ _03035_ _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09220_ _04512_ _00458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_45_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06432_ _02043_ _02059_ _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06363_ _02008_ _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09151_ net278 _04472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05314_ _00962_ _00987_ _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08102_ net587 net709 _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09082_ net152 _04416_ _04425_ _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06294_ _01916_ _01941_ _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08033_ ci_neuron.uut_simple_neuron.titan_id_1\[5\] ci_neuron.uut_simple_neuron.titan_id_0\[5\]
+ _03591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_142_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05245_ _00907_ _00920_ _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05176_ _00798_ _00818_ _00853_ _00843_ _00834_ _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_3_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09984_ _00499_ clknet_leaf_26_sys_clock_i ci_neuron.input_memory\[1\]\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08935_ net392 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08866_ internal_ih.byte1\[5\] net369 _04270_ _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07817_ net704 ci_neuron.uut_simple_neuron.titan_id_3\[29\] _03413_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08797_ _04046_ _01150_ _04231_ _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_4_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07748_ ci_neuron.uut_simple_neuron.titan_id_4\[18\] ci_neuron.uut_simple_neuron.titan_id_3\[18\]
+ _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_121_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07679_ ci_neuron.uut_simple_neuron.titan_id_4\[6\] net295 ci_neuron.uut_simple_neuron.titan_id_4\[5\]
+ ci_neuron.uut_simple_neuron.titan_id_3\[5\] _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__09521__I2 _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09418_ _03756_ net61 _00847_ _01961_ _04644_ _04645_ _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_54_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09349_ _04375_ net394 _04353_ _04588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_23_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05471__A2 _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10124_ _00248_ clknet_leaf_36_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[30\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06971__A2 _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08548__I0 _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10055_ net234 clknet_leaf_121_sys_clock_i ci_neuron.output_val_internal\[24\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08712__A3 _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08476__A2 _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06487__A1 _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold107 _04451_ net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold118 ci_neuron.uut_simple_neuron.titan_id_6\[13\] net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold129 _00284_ net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05030_ ci_neuron.address_i\[21\] ci_neuron.address_i\[20\] ci_neuron.address_i\[19\]
+ ci_neuron.address_i\[18\] _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_21_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08978__S _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06981_ _02554_ _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08539__I0 ci_neuron.value_i\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05932_ _01556_ _01591_ _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08720_ _04171_ _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05863_ _01342_ ci_neuron.uut_simple_neuron.x2\[22\] ci_neuron.uut_simple_neuron.x2\[23\]
+ _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_TAPCELL_ROW_68_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08651_ ci_neuron.uut_simple_neuron.x0\[31\] _03920_ _04114_ _04121_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07602_ _03172_ _03173_ _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05794_ _01413_ _01454_ _01455_ _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08582_ _04061_ _04062_ _04063_ _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07533_ _03100_ _03103_ _03158_ _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07464_ _03090_ _03091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08726__B _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold518_I ci_neuron.uut_simple_neuron.x0\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06415_ _02043_ _02059_ _02060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_91_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09203_ _04488_ _04503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07395_ _02557_ _02808_ _03023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09134_ _04463_ _00421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06346_ _01991_ _01969_ _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06277_ _01902_ _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_79_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09065_ _04389_ _04409_ _04410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05228_ _00833_ _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold630 ci_neuron.uut_simple_neuron.titan_id_1\[19\] net663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08461__B _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08016_ _03578_ _00151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_92_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold641 _03625_ net674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold652 _03693_ net685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_9_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold663 _03552_ net696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold685 _03378_ net718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05159_ _00837_ _00838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold674 _03323_ net707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold696 _03478_ net729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09967_ _00482_ clknet_leaf_80_sys_clock_i ci_neuron.input_memory\[1\]\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09578__S1 _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08918_ net455 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09898_ _00017_ net13 ci_neuron.address_i\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_123_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08849_ _04257_ _04264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_28_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09311__I _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05141__A1 _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_114_sys_clock_i_I clknet_4_9_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07197__A2 _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10107_ _00231_ clknet_4_15_0_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10038_ net169 clknet_leaf_77_sys_clock_i ci_neuron.output_val_internal\[7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08449__A2 _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06200_ _01836_ _01839_ _01851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_140_Right_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07180_ _02803_ _02810_ _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_42_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06131_ _01740_ _01776_ _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06062_ _01705_ _01718_ _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_14_0_sys_clock_i clknet_0_sys_clock_i clknet_4_14_0_sys_clock_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05013_ internal_ih.byte3\[5\] _00701_ _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_41_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09821_ _00400_ clknet_leaf_132_sys_clock_i internal_ih.current_instruction\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09752_ _00331_ clknet_leaf_131_sys_clock_i internal_ih.byte0\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold370_I internal_ih.byte5\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06964_ _01833_ _02535_ _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08703_ internal_ih.spi_rx_byte_i\[7\] _04148_ _04165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06895_ _01824_ _02481_ _02530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05915_ _01574_ _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09683_ _00270_ clknet_leaf_28_sys_clock_i ci_neuron.uut_simple_neuron.x3\[20\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05846_ _01445_ _01504_ _01506_ _01507_ _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_clkbuf_leaf_33_sys_clock_i_I clknet_4_4_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08634_ _03903_ _04106_ _04107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05777_ _01437_ _01439_ _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08565_ _03824_ _04043_ _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07516_ _03142_ _00247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout13 net14 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08496_ ci_neuron.value_i\[7\] _03952_ _03989_ _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xfanout24 net31 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07447_ _03001_ _03027_ _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07378_ _02863_ net447 _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06329_ _01945_ _01972_ _01975_ _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_33_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09117_ net383 _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06623__A1 _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09048_ net190 _04381_ _04394_ _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold471 internal_ih.byte0\[6\] net504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold460 internal_ih.byte2\[1\] net493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold493 internal_ih.byte0\[2\] net526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold482 internal_ih.spi_rx_byte_i\[1\] net515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_leaf_102_sys_clock_i_I clknet_4_8_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04937__A1 internal_ih.byte6\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05362__A1 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07103__A2 ci_neuron.uut_simple_neuron.x3\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09968__CLK clknet_4_12_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06680_ _02315_ _02318_ _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05700_ _01331_ _01363_ _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05631_ _01286_ _01296_ _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08350_ net745 _00182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07301_ _02927_ _02800_ _02929_ _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05562_ _01222_ _01229_ _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_47_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05493_ _01123_ _01162_ _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08281_ _03785_ _03799_ _03800_ _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08842__A2 _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07232_ _02625_ _02860_ _02861_ _02862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_4_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07163_ _02743_ _02747_ _02793_ _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06114_ _01700_ _01769_ _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_76_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07094_ _02620_ _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_clkbuf_leaf_21_sys_clock_i_I clknet_4_3_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06045_ _01665_ _01673_ _01701_ _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05959__A3 _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold585_I ci_neuron.uut_simple_neuron.titan_id_5\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08358__A1 _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07030__A1 _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09804_ _00383_ clknet_leaf_142_sys_clock_i internal_ih.byte6\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04919__B2 internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07996_ ci_neuron.uut_simple_neuron.titan_id_2\[27\] ci_neuron.uut_simple_neuron.titan_id_5\[27\]
+ ci_neuron.uut_simple_neuron.titan_id_2\[26\] ci_neuron.uut_simple_neuron.titan_id_5\[26\]
+ _03562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06947_ _02521_ _02581_ _02582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09735_ _00314_ clknet_leaf_28_sys_clock_i ci_neuron.uut_simple_neuron.x2\[16\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_65_sys_clock_i clknet_4_13_0_sys_clock_i clknet_leaf_65_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09666_ _00253_ clknet_leaf_65_sys_clock_i ci_neuron.uut_simple_neuron.x3\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06878_ _02474_ _02513_ _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_87_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08617_ _03893_ _04082_ _04092_ _03959_ _04093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_38_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05829_ _01078_ _01490_ _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09597_ net303 net122 _04790_ _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08548_ _04034_ _02335_ _04028_ _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08479_ _03957_ _03974_ _03975_ _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_118_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08597__A1 _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_131_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold290 ci_neuron.output_memory\[20\] net323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_129_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08521__A1 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09321__I0 _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08824__A2 _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08588__A1 _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09624__I1 ci_neuron.output_memory\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07850_ net591 _03438_ _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06801_ _02040_ _02437_ _02438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07781_ _03381_ _03382_ _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08760__A1 _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_107_sys_clock_i clknet_4_8_0_sys_clock_i clknet_leaf_107_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_04993_ internal_ih.byte2\[4\] _00691_ _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_39_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06732_ _02328_ _02346_ _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput3 spi_pico_i net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09520_ ci_neuron.output_memory\[22\] _04722_ _04733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06663_ _02301_ _02302_ _02303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09451_ _00727_ _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05614_ _01278_ _01280_ _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06594_ _02225_ _02234_ _02235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08402_ _03891_ _03903_ _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09382_ net213 _04611_ _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07079__A1 _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05545_ _00888_ _01142_ _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09312__I0 _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08333_ _03823_ _03835_ _03833_ _03837_ _03845_ _03846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_52_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08264_ _03771_ net124 _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05476_ _01145_ _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_144_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07215_ _02843_ _02844_ _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_132_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08195_ _00706_ _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07146_ _02775_ _02583_ _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_131_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07077_ _02656_ _02696_ _02708_ _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_112_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06028_ _01647_ _01685_ _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_58_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_4_sys_clock_i_I clknet_4_1_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_14_sys_clock_i clknet_4_1_0_sys_clock_i clknet_leaf_14_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09718_ _00297_ clknet_leaf_97_sys_clock_i internal_ih.received_byte_count\[7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07979_ net498 _03542_ net625 _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07306__A2 _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08503__A1 _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09649_ _04823_ _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_67_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_13_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06293__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09606__I1 net311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_76_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08990__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04851__I0 internal_ih.byte4\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10286_ _00579_ clknet_leaf_128_sys_clock_i ci_neuron.stream_o\[28\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09385__I3 _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07545__A2 _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08742__A1 _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09542__I0 _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_109_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_85_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05330_ _00968_ _00985_ _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_84_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07481__A1 _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05261_ _00747_ _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07000_ _02593_ _02596_ _02633_ _02634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_113_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_94_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05192_ _00835_ _00864_ _00869_ _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08951_ _04311_ _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07902_ net378 _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08882_ net334 net470 _04280_ _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_hold283_I ci_neuron.output_memory\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07833_ _03421_ _03422_ _03424_ _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold450_I ci_neuron.uut_simple_neuron.titan_id_5\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07764_ net575 ci_neuron.uut_simple_neuron.titan_id_3\[21\] _03369_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04976_ internal_ih.byte1\[5\] _00680_ _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06715_ _02351_ _02353_ _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_07695_ _03308_ _03309_ _03310_ _03311_ _03312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09503_ _04701_ _04718_ _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06646_ _02227_ ci_neuron.uut_simple_neuron.x3\[14\] ci_neuron.uut_simple_neuron.x3\[15\]
+ _02286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_84_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09434_ net111 _04655_ _04660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06577_ _01882_ _02217_ _02218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09365_ _04599_ _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05528_ _01170_ _01196_ _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09296_ _03994_ _04553_ _04558_ _00488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08316_ _03810_ _03823_ _03821_ _03831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_34_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06275__A2 _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05459_ _00961_ _01127_ _01128_ _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08247_ ci_neuron.uut_simple_neuron.x0\[9\] _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08178_ _03705_ _03710_ _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09213__A2 _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07129_ _02707_ _02709_ _02760_ _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_95_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10140_ _00205_ clknet_leaf_54_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10071_ _00198_ clknet_leaf_81_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_126_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07463__A1 _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10269_ _00562_ clknet_leaf_112_sys_clock_i ci_neuron.stream_o\[11\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05529__A1 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07480_ _02436_ _02454_ _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06500_ ci_neuron.uut_simple_neuron.x3\[11\] _02142_ _02143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_48_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06431_ _00162_ _02074_ _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06362_ _01852_ _02007_ _02008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_84_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09150_ _04471_ _00429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06293_ _01919_ _01940_ _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05313_ _00966_ _00986_ _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08101_ ci_neuron.uut_simple_neuron.titan_id_1\[16\] net708 _03649_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09081_ _04382_ _04422_ _04424_ _04411_ _04425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_05244_ _00908_ _00919_ _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08032_ net573 net688 _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05175_ _00840_ _00841_ _00852_ _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_hold498_I ci_neuron.uut_simple_neuron.x3\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09983_ _00498_ clknet_leaf_25_sys_clock_i ci_neuron.input_memory\[1\]\[18\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08934_ internal_ih.byte5\[2\] net391 _04312_ _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08865_ _04273_ _00342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07816_ net704 ci_neuron.uut_simple_neuron.titan_id_3\[29\] _03412_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08796_ _04233_ _00313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07747_ net712 _00104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04959_ _00672_ _00060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10220__D _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07678_ _03287_ _03296_ _03297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09521__I3 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06629_ _02221_ _02239_ _02269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_121_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09417_ _04606_ _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09348_ _04587_ _00511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_23_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09279_ _03955_ _04544_ _04548_ _00481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07996__A2 ci_neuron.uut_simple_neuron.titan_id_5\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10123_ _00247_ clknet_leaf_36_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08548__I1 _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10054_ net176 clknet_leaf_114_sys_clock_i ci_neuron.output_val_internal\[23\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_106_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold108 _00410_ net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07987__A2 net618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold119 ci_neuron.stream_o\[28\] net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_42_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06980_ _02560_ _02563_ _02613_ _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_95_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05931_ _01560_ _01590_ _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_13_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05862_ _01521_ _01484_ _01522_ _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08650_ _04120_ _00280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07601_ _03165_ _03171_ _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05793_ _01412_ _01438_ _01455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08581_ ci_neuron.value_i\[19\] _04032_ _04063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07532_ _03080_ _03098_ _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09874__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07463_ _03087_ _03089_ _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06414_ _02054_ _02058_ _02059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_119_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09202_ _03984_ _04494_ _04502_ _00450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_22_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07394_ _02557_ _02808_ _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09133_ net150 _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_20_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06345_ _01957_ _01991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06276_ _01921_ _01922_ _01923_ _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_79_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07978__A2 net624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09064_ ci_neuron.output_val_internal\[27\] ci_neuron.output_val_internal\[19\] ci_neuron.output_val_internal\[11\]
+ ci_neuron.output_val_internal\[3\] _04390_ _04391_ _04409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05227_ _00903_ _00227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold620 _03276_ net653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_4_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08015_ net553 net779 _03577_ _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_05158_ _00833_ _00836_ _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_92_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold642 ci_neuron.uut_simple_neuron.x2\[8\] net675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold653 ci_neuron.input_memory\[1\]\[16\] net764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold631 _03668_ net664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold675 ci_neuron.uut_simple_neuron.titan_id_0\[16\] net708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold686 ci_neuron.uut_simple_neuron.titan_id_1\[24\] net719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold664 ci_neuron.uut_simple_neuron.titan_id_1\[29\] net697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold697 internal_ih.expected_byte_count\[3\] net730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05089_ _00734_ _00765_ _00770_ _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09966_ _00481_ clknet_leaf_80_sys_clock_i ci_neuron.input_memory\[1\]\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08917_ internal_ih.byte4\[3\] net454 _04301_ _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09897_ _00012_ net13 ci_neuron.address_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08848_ _04263_ _00335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_123_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08779_ _03994_ _04218_ _04223_ _00306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_28_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_40_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_138_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09407__A2 _04636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_3_0_sys_clock_i clknet_0_sys_clock_i clknet_4_3_0_sys_clock_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07969__A2 net497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10106_ _00230_ clknet_leaf_53_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10037_ net143 clknet_leaf_77_sys_clock_i ci_neuron.output_val_internal\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06130_ _01783_ _01784_ _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06061_ _01663_ _01717_ _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05012_ _00702_ _00053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09820_ _00399_ clknet_leaf_134_sys_clock_i internal_ih.current_instruction\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09582__A1 _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06963_ _02121_ _02103_ _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09751_ _00330_ clknet_leaf_132_sys_clock_i internal_ih.byte0\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_4_0_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05914_ _01475_ _01573_ _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08702_ net130 _04136_ _04157_ internal_ih.spi_rx_byte_i\[6\] _04164_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06894_ _02074_ _02480_ _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09682_ _00269_ clknet_4_7_0_sys_clock_i ci_neuron.uut_simple_neuron.x3\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05845_ _01408_ _01503_ _01507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06699__A2 ci_neuron.uut_simple_neuron.x3\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08633_ _03900_ _04102_ _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05776_ _01389_ _01438_ _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05371__A2 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08564_ _03840_ _04044_ _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07515_ _03066_ _03141_ _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08495_ _03951_ _03987_ _03988_ _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xfanout14 net15 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout25 net26 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07446_ _03040_ _03053_ _03072_ _03073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07377_ _02868_ _02937_ _03005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_33_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06328_ _01920_ _01973_ _01974_ _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09116_ _04454_ _00412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06623__A2 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09047_ _04382_ _04388_ _04393_ _04354_ _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_32_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06259_ _01907_ _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold450 ci_neuron.uut_simple_neuron.titan_id_5\[20\] net483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold472 internal_ih.byte0\[0\] net505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_25_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold461 _04289_ net494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold483 internal_ih.byte5\[0\] net516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold494 internal_ih.byte3\[1\] net527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09949_ _00464_ clknet_leaf_18_sys_clock_i ci_neuron.uut_simple_neuron.x0\[20\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06139__A1 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_106_sys_clock_i clknet_4_8_0_sys_clock_i clknet_leaf_106_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05630_ _01261_ _01295_ _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09232__I _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07300_ _02928_ _02865_ _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05561_ _01225_ _01228_ _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06302__A1 _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05492_ _01158_ _01161_ _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_08280_ _03789_ _03792_ _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07231_ _02858_ _02859_ _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09912__CLK net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07162_ _02724_ _02742_ _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04864__A1 internal_ih.byte7\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06113_ _01749_ _01768_ _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_76_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07093_ _02680_ _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08850__I0 internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06044_ _01700_ _01675_ _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08512__S _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09803_ _00382_ clknet_leaf_141_sys_clock_i internal_ih.byte6\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_105_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07995_ _03547_ _03560_ _03545_ _03561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06946_ _02522_ _02581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_119_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09734_ _00313_ clknet_leaf_47_sys_clock_i ci_neuron.uut_simple_neuron.x2\[15\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06877_ _02512_ _02484_ _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09665_ _00252_ clknet_leaf_65_sys_clock_i ci_neuron.uut_simple_neuron.x3\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05828_ _01453_ _01489_ _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08616_ _03876_ _03879_ _04082_ _04092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_38_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09596_ _04793_ _00553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05759_ _01375_ _01337_ _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08547_ _03952_ _04031_ _04033_ _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_119_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08478_ net768 _03948_ _03975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07429_ _02920_ _02972_ _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_134_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_114_Left_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_131_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold280 internal_ih.instruction_received net313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__09546__A1 ci_neuron.output_memory\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold291 _04817_ net324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_129_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08521__A2 _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06800_ _02005_ _02436_ _02437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07780_ net445 ci_neuron.uut_simple_neuron.titan_id_3\[24\] _03382_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04992_ _00685_ _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06731_ _02316_ _02368_ _02369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09450_ _04597_ _04673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06662_ _02244_ _02255_ _02300_ _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08401_ net417 _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold159_I ci_neuron.output_val_internal\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05613_ _01240_ _01245_ _01279_ _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06593_ _02136_ _02233_ _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_4_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09381_ _04603_ _04614_ _04615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_145_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05544_ _01210_ _01211_ _01212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08332_ _03838_ _03845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout27_I net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08263_ _03784_ _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07214_ _02778_ _02841_ _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_144_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05475_ _01099_ _01102_ _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_55_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08194_ net32 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07145_ _02301_ _02307_ _02585_ _02775_ _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_113_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07076_ _02658_ _02695_ _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06027_ _01682_ _01684_ _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07978_ ci_neuron.uut_simple_neuron.titan_id_2\[24\] net624 _03547_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06929_ _02560_ _02563_ _02564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09717_ _00296_ clknet_leaf_100_sys_clock_i internal_ih.received_byte_count\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_94_sys_clock_i_I clknet_4_10_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08503__A2 _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09648_ net190 net314 _04821_ _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09579_ _04768_ _04782_ _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08814__I0 _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10285_ _00578_ clknet_leaf_129_sys_clock_i ci_neuron.stream_o\[27\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04851__I1 internal_ih.byte3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08886__I _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05260_ _00908_ _00919_ _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05191_ _00865_ net42 _00868_ _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_24_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08950_ _04321_ _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_135_Right_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07901_ _03481_ net377 _03483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09230__I0 _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08881_ _04282_ _00349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08733__A2 _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold276_I ci_neuron.output_memory\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07832_ net567 ci_neuron.uut_simple_neuron.titan_id_5\[1\] _03424_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07763_ _03364_ _03366_ _03367_ _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09502_ _03852_ ci_neuron.input_memory\[1\]\[19\] _01264_ _02552_ _04716_ _04717_
+ _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_04975_ _00681_ _00036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06714_ _02259_ _02298_ _02352_ _02353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_116_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07694_ ci_neuron.uut_simple_neuron.titan_id_4\[8\] ci_neuron.uut_simple_neuron.titan_id_3\[8\]
+ _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_84_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06645_ _02226_ _02231_ _02284_ _02285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_84_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09433_ _04652_ _04658_ _04659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09364_ _00727_ _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06576_ _01954_ _02192_ _02216_ _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__09297__I0 _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08315_ net542 _03823_ _03816_ _03818_ _03814_ _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_118_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05527_ _01172_ _01195_ _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09295_ net59 _04556_ _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05458_ _01084_ _01085_ _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08246_ _03769_ _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_133_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10218__D _00115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08177_ _03711_ _00085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07128_ _02716_ _02718_ _02759_ _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_132_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05389_ _01035_ _01057_ _01060_ _01008_ _01061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA_clkbuf_leaf_82_sys_clock_i_I clknet_4_14_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07059_ _02184_ _02691_ _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05395__I _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06983__A1 _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09221__I0 _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10070_ _00197_ clknet_leaf_80_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07932__B1 _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07463__A2 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10268_ _00561_ clknet_leaf_99_sys_clock_i ci_neuron.stream_o\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08715__A2 _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10199_ _00125_ clknet_leaf_58_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06430_ _02038_ _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06361_ _01902_ _01844_ _02007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06292_ _01920_ _01924_ _01939_ _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_05312_ _00968_ _00974_ _00985_ _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08100_ _03643_ _03645_ _03647_ _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_56_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09080_ _04389_ _04423_ _04424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05243_ _00909_ _00918_ _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08031_ net574 _00089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05174_ _00741_ _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09982_ _00497_ clknet_leaf_25_sys_clock_i ci_neuron.input_memory\[1\]\[17\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08933_ _04311_ _04312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08706__A2 _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08864_ net470 net552 _04270_ _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07815_ net705 _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08795_ _04040_ _01098_ _04231_ _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07746_ _03352_ net711 _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04958_ internal_ih.byte0\[5\] _00670_ _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_95_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_70_sys_clock_i_I clknet_4_12_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07677_ _03288_ _03293_ _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09416_ _04604_ _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_04889_ _00630_ _00012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06628_ _02266_ _02267_ _02268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_121_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06559_ _00163_ _02121_ _02153_ _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_75_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09347_ _04122_ net375 _04583_ _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_23_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09278_ net79 _04546_ _04548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08229_ ci_neuron.uut_simple_neuron.x0\[7\] _03755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10122_ _00246_ clknet_4_5_0_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_29_sys_clock_i_I clknet_4_5_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10053_ net172 clknet_leaf_120_sys_clock_i ci_neuron.output_val_internal\[22\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold109 ci_neuron.output_val_internal\[6\] net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05930_ _01563_ _01589_ _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05861_ _00780_ _01469_ _01482_ _01522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_63_sys_clock_i clknet_4_15_0_sys_clock_i clknet_leaf_63_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07600_ _03216_ _03223_ _03224_ _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_89_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08580_ _03839_ _04049_ _04026_ _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_1_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07531_ _03106_ _03116_ _03156_ _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05792_ _01421_ _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07124__A1 _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07462_ _02937_ _03088_ _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_06413_ _02057_ _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07393_ _03016_ _03020_ _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_85_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09201_ _03754_ _04500_ _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06344_ _01958_ _01968_ _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09132_ _04462_ _00420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08624__A1 _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06275_ _01899_ _01908_ _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09063_ _04383_ ci_neuron.stream_o\[3\] ci_neuron.stream_o\[19\] _04384_ _04407_
+ _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_32_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05226_ _00878_ _00882_ _00902_ _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_71_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold621 ci_neuron.uut_simple_neuron.titan_id_1\[8\] net654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold610 _03681_ net643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08014_ _03573_ net514 _03576_ _03577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05157_ ci_neuron.uut_simple_neuron.x2\[2\] ci_neuron.uut_simple_neuron.x2\[3\] ci_neuron.uut_simple_neuron.x2\[4\]
+ _00793_ _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold643 ci_neuron.uut_simple_neuron.x0\[16\] net676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold632 _03860_ net745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_12_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_92_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold676 _03649_ net709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold665 _03710_ net698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold687 _03685_ net720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__05610__A1 _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05088_ _00760_ _00767_ _00769_ _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xhold698 ci_neuron.uut_simple_neuron.titan_id_2\[6\] net731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09965_ _00480_ clknet_leaf_80_sys_clock_i ci_neuron.input_memory\[1\]\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08916_ _04302_ _00364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09896_ _00001_ net20 ci_neuron.address_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09352__A2 _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08847_ net369 net534 _04258_ _04263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_123_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08778_ _00867_ _04221_ _04223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_28_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07729_ net558 _00101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_17_sys_clock_i_I clknet_4_1_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09256__S _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10105_ _00229_ clknet_leaf_53_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_105_sys_clock_i clknet_4_8_0_sys_clock_i clknet_leaf_105_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10036_ net178 clknet_leaf_78_sys_clock_i ci_neuron.output_val_internal\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10141__D _00206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06060_ _01709_ _01716_ _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_50_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05011_ internal_ih.byte3\[4\] _00701_ _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_12_sys_clock_i clknet_4_4_0_sys_clock_i clknet_leaf_12_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06962_ net45 _02594_ _02595_ _02596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09750_ _00329_ clknet_leaf_32_sys_clock_i ci_neuron.uut_simple_neuron.x2\[31\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05913_ _01532_ _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09681_ _00268_ clknet_leaf_24_sys_clock_i ci_neuron.uut_simple_neuron.x3\[18\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08701_ _04133_ net148 _04163_ _00288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06893_ _02484_ _02512_ _02527_ _02528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08632_ _03229_ _03941_ _04105_ _00277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05844_ _01403_ _01505_ _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05775_ _00886_ _01178_ _01421_ _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08563_ _04047_ _00266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07514_ _03068_ _03140_ _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08494_ _03753_ _03976_ _03755_ _03988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07445_ _02998_ _03039_ _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout26 net27 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout15 net16 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07376_ _03002_ _03003_ _03004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_73_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06327_ _01924_ _01939_ _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09115_ net266 _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06258_ _01853_ _01906_ _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_60_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09046_ _04389_ _04392_ _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05209_ _00859_ _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06189_ _01821_ _01837_ _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold440 ci_neuron.uut_simple_neuron.titan_id_2\[13\] net473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold451 _03518_ net484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold462 internal_ih.byte3\[0\] net495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold473 ci_neuron.uut_simple_neuron.x3\[29\] net506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold495 ci_neuron.uut_simple_neuron.x0\[3\] net528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold484 _04309_ net517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09948_ _00463_ clknet_leaf_20_sys_clock_i ci_neuron.uut_simple_neuron.x0\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09879_ _00039_ net28 ci_neuron.value_i\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10019_ net78 clknet_leaf_19_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05560_ _00749_ _01227_ _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05491_ _01078_ _01159_ _01160_ _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_86_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07230_ _02858_ _02859_ _02860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07161_ _02790_ _02758_ _02791_ _02792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_125_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06112_ _01762_ _01767_ _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_140_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07092_ _02721_ _02722_ _02723_ _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_76_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06043_ _01661_ _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09555__A2 _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold473_I ci_neuron.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09802_ _00381_ clknet_leaf_137_sys_clock_i internal_ih.byte6\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07994_ ci_neuron.uut_simple_neuron.titan_id_2\[25\] ci_neuron.uut_simple_neuron.titan_id_5\[25\]
+ _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06945_ _02464_ _02463_ net47 _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07318__A1 _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09733_ _00312_ clknet_leaf_47_sys_clock_i ci_neuron.uut_simple_neuron.x2\[14\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06876_ _02487_ _02511_ _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09664_ _00251_ clknet_leaf_54_sys_clock_i ci_neuron.uut_simple_neuron.x3\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold738_I _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05827_ _01456_ _01488_ _01489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_87_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08615_ ci_neuron.value_i\[25\] _04032_ _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09595_ net98 net82 _04790_ _04793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09423__I _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05758_ _01377_ _01419_ net35 _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08546_ ci_neuron.value_i\[14\] _04032_ _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05689_ _01316_ _01317_ _01352_ _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_92_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08477_ _03971_ _03972_ _03973_ _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07428_ _02920_ _02972_ _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07359_ _02781_ _02834_ _02987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_118_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09029_ _04374_ _04376_ _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold270 ci_neuron.stream_o\[3\] net303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold281 ci_neuron.output_memory\[25\] net314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold292 ci_neuron.output_memory\[11\] net325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_129_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07309__A1 _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_58_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09537__A2 _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04991_ _00690_ _00043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06730_ _02364_ _02367_ _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_127_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06661_ _02244_ _02255_ _02300_ _02301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_78_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09243__I _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05612_ _01235_ _01239_ _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08400_ _03903_ _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06592_ _02230_ _02232_ _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_52_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09380_ _00706_ ci_neuron.input_memory\[1\]\[1\] _00745_ _01848_ _04605_ _04607_
+ _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_15_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05543_ _01011_ _01140_ _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_86_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08331_ _03836_ net390 _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_19_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05474_ _01137_ _01143_ _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_82_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08262_ _03783_ _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_52_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07213_ _02779_ _02839_ _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08193_ net163 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07144_ _02772_ _02701_ _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_07075_ _01889_ _02655_ _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06026_ _01594_ _01633_ _01683_ _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__04850__I _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07977_ net790 _03545_ _03546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06928_ _02562_ _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09716_ net211 clknet_leaf_101_sys_clock_i internal_ih.received_byte_count\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06859_ _02384_ _02448_ _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_97_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09647_ _04822_ _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09578_ ci_neuron.uut_simple_neuron.x0\[31\] ci_neuron.input_memory\[1\]\[31\] ci_neuron.uut_simple_neuron.x2\[31\]
+ ci_neuron.uut_simple_neuron.x3\[31\] _04604_ _04606_ _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_38_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08529_ _04018_ _00261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_13_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08814__I1 _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10284_ _00577_ clknet_leaf_129_sys_clock_i ci_neuron.stream_o\[26\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_144_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09542__I2 _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06269__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09207__A1 _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05492__A2 _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05190_ _00812_ _00846_ _00867_ _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_52_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_133_Left_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07900_ ci_neuron.uut_simple_neuron.titan_id_2\[12\] net376 _03482_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08880_ net269 net510 _04280_ _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07831_ net569 _00138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07762_ ci_neuron.uut_simple_neuron.titan_id_4\[20\] ci_neuron.uut_simple_neuron.titan_id_3\[20\]
+ _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09501_ _04668_ _04717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04974_ internal_ih.byte1\[4\] _00680_ _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_142_Left_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06713_ _02262_ _02297_ _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07693_ ci_neuron.uut_simple_neuron.titan_id_4\[8\] ci_neuron.uut_simple_neuron.titan_id_3\[8\]
+ net521 ci_neuron.uut_simple_neuron.titan_id_3\[7\] _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_06644_ _02227_ _02283_ _02284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_84_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09432_ _03772_ net58 _00896_ _02089_ _04644_ _04645_ _04658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_52_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06575_ _01955_ _02085_ _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05180__A1 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09363_ _04597_ _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05526_ _01183_ _01194_ _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08314_ _03829_ _00177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09294_ _03990_ _04553_ _04557_ _00487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05457_ _01084_ _01085_ _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08245_ net195 _03769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05388_ _01059_ _01060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08176_ _03709_ net698 _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09349__S _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07127_ _02720_ _02748_ _02758_ _02759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_113_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07058_ _02190_ _02690_ _02691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06009_ ci_neuron.uut_simple_neuron.x2\[28\] _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_126_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08799__I0 _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10267_ _00560_ clknet_leaf_110_sys_clock_i ci_neuron.stream_o\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_62_sys_clock_i clknet_4_14_0_sys_clock_i clknet_leaf_62_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_139_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10198_ _00124_ clknet_leaf_58_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08479__A2 _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06360_ _02005_ _01997_ _02006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06291_ _01929_ _01935_ _01938_ _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_126_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05311_ _00942_ _00984_ _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_4_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05242_ _00852_ _00912_ _00917_ _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08030_ net573 ci_neuron.uut_simple_neuron.titan_id_0\[5\] _03588_ _03589_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_142_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05173_ _00806_ _00848_ _00849_ _00829_ _00850_ _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_12_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09981_ _00496_ clknet_leaf_24_sys_clock_i ci_neuron.input_memory\[1\]\[16\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08932_ _04256_ _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_hold386_I internal_ih.byte3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04976__A1 internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08863_ net442 _00341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07814_ net704 ci_neuron.uut_simple_neuron.titan_id_3\[29\] _03410_ _03411_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08794_ _04232_ _00312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07745_ ci_neuron.uut_simple_neuron.titan_id_4\[18\] net710 _03353_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04957_ _00671_ _00059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07676_ ci_neuron.uut_simple_neuron.titan_id_4\[6\] net295 _03295_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04888_ internal_ih.byte4\[1\] _00625_ _00628_ internal_ih.byte0\[1\] _00630_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09415_ ci_neuron.output_memory\[7\] _04628_ _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06627_ _01921_ _02263_ _02264_ _02267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_121_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06558_ _02124_ _02152_ _02200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09346_ _04586_ _00510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__04900__B2 internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04900__A1 internal_ih.byte4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06489_ _02098_ _02132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05509_ _01177_ _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_90_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09277_ _03947_ _04544_ _04547_ _00480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08228_ _03753_ _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08159_ net684 net788 _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10121_ _00245_ clknet_leaf_37_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_104_sys_clock_i clknet_4_8_0_sys_clock_i clknet_leaf_104_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_100_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10052_ net189 clknet_leaf_115_sys_clock_i ci_neuron.output_val_internal\[21\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06708__A2 _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07381__A2 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10139__D _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_11_sys_clock_i clknet_4_4_0_sys_clock_i clknet_leaf_11_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__04958__A1 internal_ih.byte0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05860_ _00780_ _01469_ _01482_ _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09361__A3 _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05791_ _01415_ _01441_ _01452_ _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07530_ _03078_ _03104_ _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07461_ ci_neuron.uut_simple_neuron.x3\[27\] ci_neuron.uut_simple_neuron.x3\[28\]
+ _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06412_ _02055_ _02056_ _02057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07392_ _02812_ _03019_ _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_85_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09200_ _03979_ _04494_ _04501_ _00449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06343_ _01988_ _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09131_ net246 _04462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09770__CLK clknet_4_2_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09062_ _04405_ _04406_ _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06274_ _01898_ _01907_ _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05225_ _00879_ _00901_ _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
Xhold600 _03305_ net633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold611 _03682_ net644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08013_ net513 net802 _03576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_130_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold644 ci_neuron.uut_simple_neuron.titan_id_3\[12\] net677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05156_ _00811_ ci_neuron.uut_simple_neuron.x2\[7\] _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold622 _03607_ net655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold633 ci_neuron.uut_simple_neuron.x0\[23\] net750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_12_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08388__A1 _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold677 ci_neuron.uut_simple_neuron.titan_id_3\[18\] net710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold655 ci_neuron.uut_simple_neuron.titan_id_0\[5\] net688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold688 ci_neuron.uut_simple_neuron.titan_id_2\[18\] net721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold666 net70 net770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_05087_ _00760_ _00768_ _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold699 ci_neuron.uut_simple_neuron.x0\[15\] net732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09964_ net302 clknet_leaf_104_sys_clock_i spi_interface_cvonk.state\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08915_ net391 net443 _04301_ _04302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09895_ _00057_ net17 ci_neuron.value_i\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05175__B _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08846_ net452 _00334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_123_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05989_ _01551_ _01642_ _01643_ _01646_ _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08777_ _03990_ _04218_ _04222_ _00305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07728_ ci_neuron.uut_simple_neuron.titan_id_4\[15\] net557 _03338_ _03339_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_68_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07659_ ci_neuron.uut_simple_neuron.titan_id_4\[3\] ci_neuron.uut_simple_neuron.titan_id_3\[3\]
+ _03281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09329_ _04085_ net81 _04572_ _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10104_ _00228_ clknet_leaf_56_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10035_ net193 clknet_leaf_111_sys_clock_i ci_neuron.output_val_internal\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08606__A2 _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05010_ _00685_ _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_74_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06961_ _02540_ _02566_ _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05912_ _01528_ _01569_ _01570_ _01571_ _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_09680_ _00267_ clknet_leaf_47_sys_clock_i ci_neuron.uut_simple_neuron.x3\[17\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08917__I0 internal_ih.byte4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08700_ internal_ih.spi_rx_byte_i\[6\] _04148_ _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06892_ _02487_ _02511_ _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08631_ _04011_ _04104_ _04105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05843_ _01497_ _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05774_ _01426_ _01432_ _01436_ _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_89_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08562_ _04046_ _02384_ _04028_ _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07513_ _03135_ _03139_ _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08493_ _03753_ _03755_ _03976_ _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_07444_ _03069_ _03070_ _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout27 net30 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout16 net24 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07375_ _02942_ _02943_ _03003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06326_ _01924_ _01939_ _01973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09114_ _04453_ _00411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06257_ _01902_ _01905_ _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09045_ ci_neuron.output_val_internal\[25\] ci_neuron.output_val_internal\[17\] ci_neuron.output_val_internal\[9\]
+ ci_neuron.output_val_internal\[1\] _04390_ _04391_ _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_130_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05208_ _00841_ _00883_ _00884_ _00744_ _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_06188_ _01821_ _01837_ _01840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold441 _03486_ net474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold452 _03519_ net485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold430 _04305_ net463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold463 _04299_ net496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold474 ci_neuron.uut_simple_neuron.titan_id_4\[31\] net507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05139_ _00744_ _00784_ _00798_ _00819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xhold485 ci_neuron.uut_simple_neuron.titan_id_1\[12\] net518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold496 ci_neuron.uut_simple_neuron.x0\[27\] net529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09947_ _00462_ clknet_leaf_21_sys_clock_i ci_neuron.uut_simple_neuron.x0\[18\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08908__I0 internal_ih.byte3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09878_ _00038_ net22 ci_neuron.value_i\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08829_ _04119_ _01793_ _04246_ _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_103_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05586__A1 _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08772__A1 _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08524__A1 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10018_ net89 clknet_leaf_25_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05490_ _01081_ _01113_ _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05510__A1 _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07160_ _02720_ _02748_ _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07263__A1 _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07091_ _02678_ _02684_ _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06111_ _01615_ _01766_ _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_14_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06042_ _01698_ _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_76_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09801_ _00380_ clknet_leaf_136_sys_clock_i internal_ih.byte6\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09732_ _00311_ clknet_leaf_47_sys_clock_i ci_neuron.uut_simple_neuron.x2\[13\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07993_ _03546_ _03558_ _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06944_ _02411_ _02356_ _02410_ _02406_ _02467_ _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__08515__A1 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06875_ _02510_ _02491_ _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09663_ _00250_ clknet_leaf_62_sys_clock_i ci_neuron.uut_simple_neuron.x3\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05826_ _01460_ _01487_ _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_87_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08614_ _04090_ _00274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_19_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09594_ net285 _00552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08545_ _04000_ _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_38_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05757_ _01104_ _01188_ _01370_ _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_05688_ _01316_ _01317_ _01352_ _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08476_ ci_neuron.value_i\[4\] _03951_ _03973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09491__A2 _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07427_ _03054_ _02996_ _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_107_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09618__I1 ci_neuron.output_memory\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07358_ _02784_ _02833_ _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_118_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06309_ _01954_ _01955_ _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_28_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10237__D _00133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07289_ _02899_ _02907_ _02917_ _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_131_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_131_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09028_ _04191_ _04375_ _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold271 ci_neuron.uut_simple_neuron.titan_id_5\[8\] net304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold260 internal_ih.received_byte_count\[2\] net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold282 ci_neuron.output_memory\[27\] net315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold293 _04804_ net326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07309__A2 ci_neuron.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09554__I0 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_142_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09306__I0 _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07493__A1 _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09609__I1 ci_neuron.output_memory\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_78_sys_clock_i_I clknet_4_11_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_46_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06599__A3 _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04990_ internal_ih.byte2\[3\] _00686_ _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06660_ _02258_ _02299_ _02300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_05611_ _01248_ _01277_ _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_35_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06591_ _02231_ net500 _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_35_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05542_ _01018_ _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08330_ _03843_ _00179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05473_ _00864_ _01142_ _01143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08261_ ci_neuron.uut_simple_neuron.x0\[11\] _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07212_ _02842_ _00243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08192_ net288 _00066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07143_ _02771_ _02768_ net39 _02704_ _02773_ _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_42_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07074_ _02706_ _00241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_125_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06025_ _01601_ _01632_ _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_100_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_89_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07976_ net789 net823 _03545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06927_ _02279_ _02561_ _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09715_ _00294_ clknet_leaf_97_sys_clock_i internal_ih.received_byte_count\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09646_ net206 net322 _04821_ _04822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06858_ _02447_ _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06789_ _01991_ _02375_ _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05809_ _00852_ _01469_ _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09577_ ci_neuron.output_memory\[31\] _04766_ _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08528_ _04017_ _02139_ _03969_ _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_136_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07475__A1 _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08459_ net32 ci_neuron.uut_simple_neuron.x0\[1\] net163 _03958_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_92_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05789__A1 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09519__A3 _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10283_ _00576_ clknet_leaf_130_sys_clock_i ci_neuron.stream_o\[25\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_61_sys_clock_i clknet_4_14_0_sys_clock_i clknet_leaf_61_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_144_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07950__A2 net414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_66_sys_clock_i_I clknet_4_13_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09542__I3 _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_54_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_135_sys_clock_i_I clknet_4_2_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07830_ _03421_ _03422_ _03423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07761_ ci_neuron.uut_simple_neuron.titan_id_4\[20\] ci_neuron.uut_simple_neuron.titan_id_3\[20\]
+ _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07941__A2 ci_neuron.uut_simple_neuron.titan_id_5\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06712_ _02350_ _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09500_ _04666_ _04716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_04973_ _00664_ _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07692_ _03300_ _03305_ _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09877__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06643_ ci_neuron.uut_simple_neuron.x3\[14\] _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09431_ ci_neuron.output_memory\[9\] _04650_ _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06574_ _02177_ _02196_ _02214_ _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09362_ _04596_ _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05525_ _01171_ _01193_ _01194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08313_ _03822_ _03824_ _03828_ _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_145_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09293_ net61 _04556_ _04557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05456_ _01082_ _01112_ _01125_ _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_74_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08244_ _03768_ _00198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05387_ _01058_ _01056_ _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08175_ net697 ci_neuron.uut_simple_neuron.titan_id_0\[29\] _03710_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_42_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07126_ _02751_ _02757_ _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_42_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07057_ _02329_ _02628_ _02689_ _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_88_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_103_sys_clock_i clknet_4_8_0_sys_clock_i clknet_leaf_103_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_101_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06008_ _01621_ _01622_ _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_126_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07959_ net524 net458 _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_98_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09629_ net380 _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_54_sys_clock_i_I clknet_4_15_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_10_sys_clock_i clknet_4_4_0_sys_clock_i clknet_leaf_10_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_55_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10266_ _00559_ clknet_leaf_112_sys_clock_i ci_neuron.stream_o\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10197_ _00123_ clknet_leaf_58_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07439__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10107__CLK clknet_4_15_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06290_ _01937_ _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05310_ _00868_ _00983_ _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_123_sys_clock_i_I clknet_4_3_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05241_ _00913_ _00916_ _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05172_ _00831_ _00844_ _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_29_sys_clock_i clknet_4_5_0_sys_clock_i clknet_leaf_29_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_3_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07611__A1 _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09980_ _00495_ clknet_leaf_23_sys_clock_i ci_neuron.input_memory\[1\]\[15\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08931_ _04310_ _00371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08862_ internal_ih.byte1\[3\] net441 _04270_ _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07813_ _03387_ _03388_ _03404_ _03409_ _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_08793_ _04034_ net755 _04231_ _04232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07744_ _03350_ _03351_ _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04956_ internal_ih.byte0\[4\] _00670_ _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07675_ net297 _00122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06626_ _02265_ _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_04887_ _00629_ _00001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09414_ _04627_ _04639_ _04641_ _04642_ _00522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_137_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09419__A2 _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06557_ _02170_ _02198_ _02199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_75_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09345_ _04119_ net338 _04583_ _04586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06488_ _02088_ _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05508_ _01173_ _01176_ _01042_ _01177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06102__A1 _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09276_ net86 _04546_ _04547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05439_ _01049_ _01050_ _01048_ _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08227_ _03752_ _03753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08158_ net684 net788 _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07109_ _02441_ _02740_ _02741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08089_ net519 _03636_ _03638_ _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_30_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10120_ _00244_ clknet_leaf_38_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[26\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10051_ net167 clknet_leaf_121_sys_clock_i ci_neuron.output_val_internal\[20\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05916__A1 _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_42_sys_clock_i_I clknet_4_7_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05080__A1 _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10249_ _00146_ clknet_leaf_16_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05907__A1 _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05790_ _01418_ _01440_ _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_4_13_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_111_sys_clock_i_I clknet_4_10_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06580__A1 _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09532__I _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07460_ _03085_ _03086_ _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_76_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06411_ _01860_ _01931_ _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07391_ _03017_ _03018_ _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09915__CLK net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06342_ _01953_ _01988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09130_ _04461_ _00419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_20_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09061_ _04358_ ci_neuron.stream_o\[11\] _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06273_ _01894_ _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08012_ _03575_ _00150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05224_ _00885_ _00900_ _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold601 _03306_ net634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold612 ci_neuron.uut_simple_neuron.titan_id_2\[16\] net645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_4_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold645 _03327_ net678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05155_ _00832_ _00833_ _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold634 ci_neuron.uut_simple_neuron.titan_id_5\[10\] net667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_69_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold623 _03608_ net656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold678 _03353_ net711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05086_ _00766_ _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold667 ci_neuron.input_memory\[1\]\[19\] net774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold656 _03593_ net689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09963_ net250 clknet_leaf_103_sys_clock_i spi_interface_cvonk.state\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold689 _03509_ net722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08914_ _04290_ _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_85_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09894_ _00056_ net17 ci_neuron.value_i\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08845_ internal_ih.byte0\[4\] net451 _04258_ _04262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08776_ _00847_ _04221_ _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08560__A2 _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05988_ _01644_ _01645_ _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07727_ _03334_ _03335_ _03337_ _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__09442__I _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04939_ internal_ih.byte6\[5\] _00658_ _00659_ internal_ih.byte2\[5\] _00661_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07658_ net716 _00118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07589_ _03145_ _03214_ _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_138_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06609_ _02209_ _02249_ _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_95_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09328_ _04079_ _04546_ _04576_ _00502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_4_11_0_sys_clock_i clknet_0_sys_clock_i clknet_4_11_0_sys_clock_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_48_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09259_ _04383_ _04373_ _04374_ _04533_ _00476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08871__I0 internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05210__I _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_30_sys_clock_i_I clknet_4_4_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10103_ _00169_ clknet_leaf_56_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09328__A1 _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10034_ net123 clknet_leaf_94_sys_clock_i ci_neuron.output_val_internal\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08862__I0 internal_ih.byte1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09406__I2 _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09567__A1 net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09527__I _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06960_ _02540_ _02566_ _02594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06891_ _02476_ _02483_ _02525_ _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05911_ _01527_ _01536_ _01571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05842_ _01408_ _01503_ _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08630_ _04101_ _04103_ _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_89_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05773_ _01425_ _01435_ _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08561_ _03996_ _04042_ _04044_ _04045_ _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_07512_ _03137_ _03138_ _03139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08492_ _03940_ _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07443_ _03041_ _03052_ _03070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06856__A2 _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout28 net30 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout17 net18 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07374_ _02932_ _02941_ _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09113_ net194 _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06325_ _01947_ _01971_ _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_33_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06256_ _01873_ _01904_ _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09044_ internal_ih.data_pointer\[1\] _04391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05207_ _00842_ _00871_ _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_hold780_I _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold420 ci_neuron.uut_simple_neuron.x0\[26\] net453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06187_ _01837_ _01838_ _01839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold453 internal_ih.spi_rx_byte_i\[3\] net486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold442 internal_ih.byte1\[5\] net475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold431 internal_ih.spi_rx_byte_i\[6\] net464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold475 _03419_ net508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05138_ _00814_ _00817_ _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold464 ci_neuron.uut_simple_neuron.titan_id_5\[23\] net497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold486 _03634_ net519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06792__A1 _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05069_ ci_neuron.uut_simple_neuron.x2\[2\] _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09946_ _00461_ clknet_leaf_21_sys_clock_i ci_neuron.uut_simple_neuron.x0\[17\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold497 internal_ih.current_instruction\[3\] net530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09877_ _00037_ net28 ci_neuron.value_i\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06544__A1 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08828_ _04251_ _00327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08759_ _00737_ _04211_ _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_103_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09283__S _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10017_ net71 clknet_leaf_22_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04954__I _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07090_ _02686_ _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06110_ _01613_ _01765_ _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06041_ _01255_ _01697_ _01698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_76_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09800_ _00379_ clknet_leaf_145_sys_clock_i internal_ih.byte6\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07992_ _03552_ _03554_ _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06943_ _02577_ _02521_ _02578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09731_ _00310_ clknet_leaf_49_sys_clock_i ci_neuron.uut_simple_neuron.x2\[12\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07971__B1 _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06874_ _02509_ _02493_ _02510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_hold459_I internal_ih.byte3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09662_ _04830_ _00582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05825_ _01467_ _01486_ _01487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08613_ _04089_ _02865_ _04086_ _04090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09593_ ci_neuron.stream_o\[1\] net284 _04790_ _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05756_ _01333_ _01372_ _01145_ _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_08544_ _03808_ _04030_ _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_38_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05687_ _01236_ _01351_ _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08475_ _03739_ _03963_ _03972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07426_ _03053_ _03040_ _03054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_135_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09079__I0 ci_neuron.output_val_internal\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07357_ _02985_ _00245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_118_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06308_ _01933_ _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07288_ _02902_ _02906_ _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_131_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09027_ _04152_ _04172_ _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06239_ _01888_ _00166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold250 internal_ih.current_instruction\[7\] net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold261 _00292_ net294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_leaf_60_sys_clock_i clknet_4_15_0_sys_clock_i clknet_leaf_60_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold272 _03464_ net305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__05017__A1 internal_ih.byte3\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold294 ci_neuron.output_memory\[30\] net327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold283 ci_neuron.output_memory\[6\] net316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_130_Right_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09929_ _00444_ clknet_leaf_77_sys_clock_i ci_neuron.uut_simple_neuron.x0\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_129_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08690__A1 _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_1_sys_clock_i_I clknet_4_1_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09490__I0 _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_79_sys_clock_i clknet_4_14_0_sys_clock_i clknet_leaf_79_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_71_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05610_ _01124_ _01276_ _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06590_ _02227_ ci_neuron.uut_simple_neuron.x3\[14\] _02231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_87_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05541_ _01180_ _01208_ _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05472_ _01139_ _01141_ _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08260_ _03776_ _03782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07211_ _02778_ _02841_ _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_144_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08808__I0 _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08191_ ci_neuron.uut_simple_neuron.titan_id_1\[2\] net287 _03723_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07142_ _02647_ _02765_ _02764_ _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_82_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07236__A2 _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07073_ _02700_ _02705_ _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06024_ _01648_ _01681_ _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09233__I0 _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_102_sys_clock_i clknet_4_8_0_sys_clock_i clknet_leaf_102_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_140_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07975_ net789 ci_neuron.uut_simple_neuron.titan_id_5\[25\] _03544_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06926_ _02232_ _02386_ _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_93_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09714_ net273 clknet_leaf_101_sys_clock_i internal_ih.received_byte_count\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06857_ _02452_ _02455_ _02492_ _02493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07235__I ci_neuron.uut_simple_neuron.x3\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09645_ _04810_ _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05808_ _01432_ _01436_ _01468_ _01469_ _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_06788_ _01969_ _02374_ _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09450__I _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09576_ _04765_ _04777_ _04779_ _04780_ _00546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05739_ _01356_ _01402_ _01354_ _01403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08527_ _04013_ _04014_ _04015_ _04016_ _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_08458_ _03940_ _03957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07409_ _03034_ _03036_ _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_135_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08389_ _03886_ _03887_ _03895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09224__I0 _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10282_ _00575_ clknet_leaf_130_sys_clock_i ci_neuron.stream_o\[24\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06910__A1 _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04921__B1 _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_139_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08415__A1 _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_28_sys_clock_i clknet_4_7_0_sys_clock_i clknet_leaf_28_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_45_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09215__I0 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07760_ net658 _00106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04972_ _00679_ _00035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06711_ _02266_ _02311_ _02349_ _02350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_79_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07691_ _03287_ _03296_ _03307_ _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_79_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09430_ _04649_ _04651_ _04654_ _04656_ _00524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06642_ _02136_ _02233_ _02281_ _02282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_94_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06573_ _02180_ _02195_ _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09361_ _04595_ _00724_ _03923_ _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_129_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05524_ _01147_ _01188_ _01189_ _01192_ _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_09292_ _04545_ _04556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08312_ _03826_ _03827_ _03828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08243_ _03766_ _03767_ _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_fanout25_I net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05455_ net41 _01111_ _01125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05386_ _00741_ _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08174_ _03704_ net681 _03708_ _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07125_ _02754_ _02756_ _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_141_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07056_ _02330_ _02494_ _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_70_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06007_ _01662_ _01664_ _01665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09445__I _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09382__A2 _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07958_ _03520_ _03525_ _03526_ _03528_ _03529_ _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_06909_ _02131_ _02543_ _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07889_ _03467_ _03468_ _03469_ _03471_ _03472_ _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_09628_ net379 ci_neuron.output_memory\[16\] _04811_ _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09559_ _00727_ _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05459__A1 _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_137_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06959__A1 _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10265_ _00558_ clknet_leaf_98_sys_clock_i ci_neuron.stream_o\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10196_ _00122_ clknet_leaf_58_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05240_ _00914_ _00915_ _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05171_ _00831_ _00844_ _00849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_141_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06889__I _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05622__A1 _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08930_ net403 net491 _04306_ _04310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08861_ _04271_ _00340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07812_ net600 ci_neuron.uut_simple_neuron.titan_id_3\[28\] _03403_ _03406_ _03408_
+ _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08792_ _04224_ _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_hold274_I ci_neuron.output_memory\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07743_ _03347_ _03348_ _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04955_ _00664_ _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07674_ _03292_ net296 _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04886_ internal_ih.byte4\[0\] _00625_ _00628_ internal_ih.byte0\[0\] _00629_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06625_ _02263_ _02264_ _01921_ _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09413_ net142 _04633_ _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_121_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06556_ _02172_ _02197_ _02198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09344_ _04585_ _00509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_23_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06487_ _01850_ _02129_ _02130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05507_ _01140_ _00981_ _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
X_09275_ _04545_ _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05438_ _01049_ _01048_ _01050_ _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_90_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08226_ ci_neuron.uut_simple_neuron.x0\[6\] _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05861__A1 _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08157_ _03694_ _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07108_ _02390_ _02615_ _02740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05369_ _01013_ _01014_ _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_73_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08088_ ci_neuron.uut_simple_neuron.titan_id_1\[13\] ci_neuron.uut_simple_neuron.titan_id_0\[13\]
+ _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07039_ _02619_ _02627_ _02672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10050_ net137 clknet_leaf_114_sys_clock_i ci_neuron.output_val_internal\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_82_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_3_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09291__A1 _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_91_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10248_ _00145_ clknet_leaf_16_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[26\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10179_ _00076_ clknet_leaf_18_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06410_ _01858_ _02055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_4_0_0_sys_clock_i clknet_0_sys_clock_i clknet_4_0_0_sys_clock_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07390_ _02676_ _02858_ _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_85_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06341_ _01985_ _01986_ _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09282__A1 _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06272_ _01891_ _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06096__A1 _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09060_ _04360_ _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05223_ _00889_ _00899_ _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08011_ _03573_ net514 _03575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold602 ci_neuron.uut_simple_neuron.titan_id_4\[4\] net635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold624 ci_neuron.uut_simple_neuron.titan_id_4\[20\] net657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_102_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05154_ ci_neuron.uut_simple_neuron.x2\[2\] ci_neuron.uut_simple_neuron.x2\[3\] ci_neuron.uut_simple_neuron.x2\[4\]
+ ci_neuron.uut_simple_neuron.x2\[5\] _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
Xhold613 _03498_ net646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold635 ci_neuron.input_memory\[1\]\[17\] net753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_69_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold679 _03354_ net712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold646 _03328_ net679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05085_ _00756_ _00766_ _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold668 ci_neuron.uut_simple_neuron.titan_id_1\[14\] net701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold657 _03595_ net690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09962_ net405 clknet_leaf_104_sys_clock_i spi_interface_cvonk.state\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_139_Left_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08913_ _04300_ _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09893_ _00054_ net23 ci_neuron.value_i\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08844_ _04261_ _00333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09870__D _00061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05987_ _01634_ _01636_ _01638_ _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_109_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08775_ _04210_ _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07726_ ci_neuron.uut_simple_neuron.titan_id_4\[14\] ci_neuron.uut_simple_neuron.titan_id_3\[14\]
+ _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_0_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04938_ _00660_ _00013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_28_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07657_ ci_neuron.uut_simple_neuron.titan_id_4\[3\] ci_neuron.uut_simple_neuron.titan_id_3\[3\]
+ net715 _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_04869_ _00605_ _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07588_ _03146_ _03213_ _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06608_ _02244_ _02248_ _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09648__I0 net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06539_ _02141_ _02181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09327_ net67 _04556_ _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09258_ _04381_ _04384_ _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08209_ _03733_ _03737_ _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09189_ _04488_ _04494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08802__I _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10102_ _00168_ clknet_leaf_56_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09328__A2 _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06322__I _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10033_ net83 clknet_leaf_94_sys_clock_i ci_neuron.output_val_internal\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_144_Right_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09406__I3 _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06890_ _02479_ _02482_ _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05910_ _01530_ _01534_ _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05841_ _01450_ _01443_ _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06553__A2 _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05772_ _01430_ _01434_ _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_77_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08560_ ci_neuron.value_i\[16\] _04001_ _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07511_ _02993_ _03055_ _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08491_ _03957_ _03984_ _03985_ _00256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07442_ _03042_ _03043_ _03051_ _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout29 net30 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout18 net23 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07373_ _02945_ _02948_ _03000_ _03001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06324_ _01951_ _01970_ _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_84_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09112_ _04415_ net140 _04452_ _00410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_33_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06255_ ci_neuron.uut_simple_neuron.x3\[5\] _01903_ _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09043_ internal_ih.data_pointer\[0\] _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_130_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06186_ ci_neuron.uut_simple_neuron.x3\[3\] _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05206_ _00853_ _00871_ _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold410 internal_ih.byte3\[2\] net443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05137_ _00781_ _00816_ _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold432 _04265_ net465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold421 internal_ih.byte3\[3\] net454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold443 internal_ih.byte1\[0\] net476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold454 ci_neuron.uut_simple_neuron.titan_id_1\[30\] net487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06241__A1 _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07238__I ci_neuron.uut_simple_neuron.x3\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold487 _03637_ net520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold476 internal_ih.byte1\[7\] net509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold465 _03541_ net498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05068_ _00737_ _00751_ _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold498 ci_neuron.uut_simple_neuron.x3\[30\] net531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09945_ _00460_ clknet_leaf_119_sys_clock_i ci_neuron.uut_simple_neuron.x0\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09876_ _00036_ net20 ci_neuron.value_i\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08827_ _04116_ net758 _04246_ _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08758_ _04210_ _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_103_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07709_ net707 _00097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08689_ net486 _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_138_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08541__I0 _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_78_sys_clock_i clknet_4_11_0_sys_clock_i clknet_leaf_78_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_101_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05035__A2 _00718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10016_ net73 clknet_leaf_23_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09363__I _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04849__A2 _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09237__A1 _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06040_ _01179_ _01696_ _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_76_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_101_sys_clock_i clknet_4_8_0_sys_clock_i clknet_leaf_101_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09538__I _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07991_ _03557_ _00146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06942_ _02463_ _02465_ _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09730_ _00309_ clknet_leaf_69_sys_clock_i ci_neuron.uut_simple_neuron.x2\[11\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09273__I _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06873_ _02505_ _02508_ _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_119_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09661_ net139 net361 _04826_ _04830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05824_ _01470_ _01485_ _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08612_ ci_neuron.value_i\[24\] _04088_ _03953_ _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09592_ net363 _00551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05755_ _01416_ _01387_ _01417_ _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08543_ _03794_ _03796_ _04015_ _04030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_38_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05337__I0 _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05686_ _01319_ _01350_ _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_106_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08474_ _03942_ _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_18_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07425_ _03041_ _03052_ _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07356_ _02979_ _02984_ _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_118_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07287_ _02910_ _02912_ _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06307_ _01931_ _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_131_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06238_ _01885_ _01887_ _01888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09026_ _04145_ _04179_ _04373_ _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06169_ _01820_ _01822_ _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold262 ci_neuron.uut_simple_neuron.titan_id_3\[6\] net295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold240 _00293_ net273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold251 ci_neuron.output_memory\[1\] net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06214__A1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold273 _03466_ net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold295 ci_neuron.output_memory\[26\] net328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold284 _04798_ net317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09928_ net222 clknet_leaf_102_sys_clock_i internal_ih.received_byte_count\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09183__I _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09554__I2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09859_ _00438_ clknet_leaf_16_sys_clock_i ci_neuron.output_memory\[27\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_142_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08690__A2 _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_27_sys_clock_i clknet_4_6_0_sys_clock_i clknet_leaf_27_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_52_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08262__I _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_91_sys_clock_i_I clknet_4_11_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05540_ _00961_ _01207_ _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05471_ _00982_ _01017_ _01140_ _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_74_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07210_ _02840_ _02841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_129_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08190_ _03722_ _00087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07141_ _02764_ _02700_ _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07072_ _02587_ _02701_ _02704_ _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_113_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06023_ _01652_ _01680_ _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06747__A2 _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold471_I internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07516__I _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07974_ _03543_ _00143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06925_ _02550_ _02559_ _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09536__I2 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09713_ net294 clknet_leaf_101_sys_clock_i internal_ih.received_byte_count\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06856_ _02444_ _02451_ _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_hold736_I _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09644_ net321 _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05807_ _01435_ _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06787_ _02369_ _02399_ _02423_ _02424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09575_ net258 _04771_ _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05738_ _01353_ _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_93_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08526_ ci_neuron.value_i\[11\] _03965_ _04016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05669_ ci_neuron.uut_simple_neuron.x2\[19\] ci_neuron.uut_simple_neuron.x2\[20\]
+ _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08457_ _03941_ _03955_ _03956_ _00251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_119_sys_clock_i_I clknet_4_3_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07408_ _02041_ _03035_ _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08388_ _03893_ _03889_ _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07339_ _01929_ _02420_ _02317_ _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06435__A1 _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05238__A2 _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09224__I1 _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09009_ internal_ih.data_pointer\[1\] _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10281_ _00574_ clknet_leaf_129_sys_clock_i ci_neuron.stream_o\[23\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06330__I _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06910__A2 _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04921__B2 internal_ih.byte1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08415__A2 _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06977__A2 _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09215__I1 _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_102_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08720__I _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06240__I _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04971_ internal_ih.byte1\[3\] _00675_ _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06710_ _02319_ _02348_ _02349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_clkbuf_leaf_38_sys_clock_i_I clknet_4_5_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07690_ _03295_ _03298_ _03307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06641_ _02279_ _02280_ _02281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_87_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06572_ _01827_ _02212_ _02213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09360_ _00708_ _00729_ _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_111_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05523_ _01190_ _01191_ _01186_ _01192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_74_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09291_ _03984_ _04553_ _04555_ _00486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08311_ _03814_ _03819_ _03827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05454_ _00934_ _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08242_ _03765_ _03761_ _03764_ _03767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_145_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout18_I net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05385_ _01056_ _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08173_ _03707_ _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07124_ _01882_ _02755_ _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08831__S _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07055_ _02687_ _02675_ _02688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_120_Left_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06006_ _01663_ _01624_ _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_107_sys_clock_i_I clknet_4_8_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08590__A1 _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07957_ ci_neuron.uut_simple_neuron.titan_id_2\[21\] net414 _03529_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_126_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06908_ _02098_ _02542_ _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07888_ ci_neuron.uut_simple_neuron.titan_id_2\[9\] ci_neuron.uut_simple_neuron.titan_id_5\[9\]
+ _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06839_ _01984_ _02009_ _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09627_ _04810_ _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_108_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09558_ _04696_ _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08509_ _04000_ _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_136_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09489_ ci_neuron.output_memory\[17\] _04698_ _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_136_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08805__I _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08540__I _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10264_ _00557_ clknet_leaf_98_sys_clock_i ci_neuron.stream_o\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10195_ _00121_ clknet_leaf_60_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08956__I0 internal_ih.byte6\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09371__I _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05404__I _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08636__A2 _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05170_ _00814_ _00847_ _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_25_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07072__A1 _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_26_sys_clock_i_I clknet_4_6_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08860_ net481 net526 _04270_ _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07811_ _03407_ _03408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08791_ _04230_ _00311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07742_ ci_neuron.uut_simple_neuron.titan_id_4\[17\] ci_neuron.uut_simple_neuron.titan_id_3\[17\]
+ _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_04954_ _00669_ _00058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07673_ ci_neuron.uut_simple_neuron.titan_id_4\[6\] net295 _03293_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05138__A1 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04885_ _00627_ _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06624_ _01871_ _02218_ _02264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09412_ _04630_ _04640_ _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_121_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09343_ _04116_ net95 _04583_ _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06555_ _02177_ _02196_ _02197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_74_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08627__A2 _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06486_ _02125_ _02128_ _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05506_ _00887_ _01142_ _01174_ _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_75_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09274_ _04542_ _04545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05437_ _01088_ _01095_ _01107_ _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08225_ net512 _00196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05368_ _01013_ _01014_ _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08156_ _03692_ net685 _03694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_132_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07107_ _02738_ _02729_ _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_28_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09669__CLK clknet_4_13_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05299_ _00971_ _00972_ _00965_ _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08087_ net520 _00068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07038_ net52 _02669_ _02670_ _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05377__A1 _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08989_ net263 _04341_ _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09418__I1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10247_ _00144_ clknet_leaf_17_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08554__A1 _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10178_ _00075_ clknet_leaf_21_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_14_sys_clock_i_I clknet_4_1_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05540__A1 _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09657__I1 net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06340_ _01830_ _01877_ _01892_ _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06271_ _01890_ _01917_ _01918_ _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06096__A2 _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05222_ _00890_ _00898_ _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_60_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08010_ net513 ci_neuron.uut_simple_neuron.titan_id_5\[30\] _03574_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold603 _03284_ net636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold625 _03365_ net658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05153_ _00787_ _00816_ _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_69_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold636 _03475_ net669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold614 net819 net647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05084_ ci_neuron.uut_simple_neuron.x2\[4\] _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold669 _03640_ net702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold658 ci_neuron.uut_simple_neuron.titan_id_1\[22\] net691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_leaf_9_sys_clock_i_I clknet_4_4_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold647 ci_neuron.uut_simple_neuron.titan_id_1\[28\] net680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09961_ net734 clknet_leaf_109_sys_clock_i internal_ih.data_pointer\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08912_ net491 net527 _04296_ _04300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09593__I0 ci_neuron.stream_o\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09892_ _00053_ net17 ci_neuron.value_i\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08843_ net441 _04155_ _04258_ _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05986_ _01634_ _01636_ _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08774_ _03984_ _04218_ _04220_ _00304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07725_ net639 _00100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09345__I0 _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04937_ internal_ih.byte6\[4\] _00658_ _00659_ internal_ih.byte2\[4\] _00660_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_28_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06859__A1 _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06323__A3 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ _03275_ _03277_ _03278_ _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04868_ _00615_ _00028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07587_ _03150_ _03212_ _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06607_ _02246_ _02247_ _02248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06538_ _02147_ _02149_ _02179_ _02180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09326_ _04575_ _00501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09257_ _04532_ _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06469_ _02030_ _02016_ _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_106_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08208_ _03734_ _03735_ _03736_ _03737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_134_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09025__A2 _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09188_ _03955_ _04489_ _04493_ _00445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08139_ _03676_ _03678_ _03679_ _03680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xclkbuf_leaf_77_sys_clock_i clknet_4_10_0_sys_clock_i clknet_leaf_77_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_105_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05598__A1 _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08784__A1 _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10101_ _00167_ clknet_leaf_55_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10032_ net214 clknet_leaf_93_sys_clock_i ci_neuron.output_val_internal\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07434__I _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09336__I0 _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09834__CLK clknet_4_11_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09297__S _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_100_sys_clock_i clknet_4_8_0_sys_clock_i clknet_leaf_100_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09016__A2 ci_neuron.stream_o\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05589__A1 _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08527__A1 _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05840_ _01307_ _01312_ _01501_ _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07510_ _03136_ _03054_ _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05771_ _01433_ _01380_ _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08490_ _01959_ _03980_ _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07441_ _03067_ _03058_ _03068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05513__A1 _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout19 net21 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07372_ _02999_ _02944_ _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06323_ _01953_ _01958_ _01969_ _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09111_ internal_ih.spi_tx_byte_o\[7\] _04427_ _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_33_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06254_ ci_neuron.uut_simple_neuron.x3\[6\] _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_119_sys_clock_i clknet_4_3_0_sys_clock_i clknet_leaf_119_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09042_ _04355_ _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06185_ ci_neuron.uut_simple_neuron.x3\[2\] _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05205_ _00879_ _00873_ _00881_ _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold411 internal_ih.byte6\[3\] net444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold400 _04292_ net433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05136_ _00794_ _00796_ _00815_ _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xhold422 _04303_ net455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_4_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold444 _04278_ net477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_25_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold433 internal_ih.byte2\[6\] net466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_40_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold477 internal_ih.byte1\[3\] net510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold466 ci_neuron.output_memory\[28\] net627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold455 _03718_ net488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold499 ci_neuron.uut_simple_neuron.titan_id_4\[19\] net532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_111_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold488 ci_neuron.uut_simple_neuron.titan_id_4\[7\] net521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05067_ _00750_ _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09944_ _00459_ clknet_leaf_118_sys_clock_i ci_neuron.uut_simple_neuron.x0\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05044__A3 _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09875_ _00035_ net28 ci_neuron.value_i\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08826_ _04250_ _00326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09191__A1 _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09318__I0 _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05969_ _01609_ _01627_ _01628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08757_ _04207_ _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_68_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07708_ net706 ci_neuron.uut_simple_neuron.titan_id_3\[11\] _03322_ _03323_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_68_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08688_ net117 _04137_ _04142_ _04152_ _04154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07639_ _03187_ _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05504__A1 _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08541__I1 _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07257__A1 _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09309_ _04565_ _00494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_26_sys_clock_i clknet_4_6_0_sys_clock_i clknet_leaf_26_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_106_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04866__I0 internal_ih.byte4\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_6_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10015_ net87 clknet_leaf_23_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09237__A2 _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07990_ net619 _03556_ _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06941_ _02573_ _02575_ _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__07971__A2 net497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09660_ _04829_ _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07074__I _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06872_ _02507_ _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_66_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08611_ _03877_ _03869_ _04077_ _04088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05734__A1 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05823_ _01471_ _01482_ _01484_ _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09591_ ci_neuron.stream_o\[0\] net362 _04790_ _04791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05754_ _01388_ _01392_ _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08542_ _04029_ _00263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08473_ _03970_ _00253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07424_ _03044_ _03051_ _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05685_ _01284_ _01349_ _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08834__S _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07355_ _02778_ _02980_ _02983_ _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_135_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06306_ _01834_ _01952_ _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07286_ _02915_ _00244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06237_ _01857_ _01864_ _01886_ _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09025_ _04178_ _00600_ _04186_ _04373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_131_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08739__A1 _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06168_ _01821_ _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold241 ci_neuron.input_memory\[1\]\[22\] net568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_13_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold230 internal_ih.current_instruction\[2\] net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold252 _04792_ net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold263 _03293_ net296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05119_ _00786_ _00789_ _00799_ _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06099_ _01754_ _01667_ ci_neuron.uut_simple_neuron.x2\[30\] _01755_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xhold285 ci_neuron.uut_simple_neuron.x0\[7\] net596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold296 ci_neuron.uut_simple_neuron.x0\[25\] net329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold274 ci_neuron.output_memory\[5\] net307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07962__A2 net458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09927_ _00032_ net5 ci_neuron.instruction_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_129_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09554__I3 _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09858_ _00437_ clknet_leaf_125_sys_clock_i ci_neuron.output_memory\[26\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08809_ _04241_ _00318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09789_ _00368_ clknet_leaf_144_sys_clock_i internal_ih.byte4\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_142_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09467__A2 _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09490__I2 _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07402__A1 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07953__A2 net414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05407__I _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05192__A2 _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05470_ _01091_ _01099_ _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_15_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07140_ _02647_ _02765_ _02764_ _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_144_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08453__I _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07071_ _02637_ _02702_ net48 _02703_ _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_140_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06022_ _01650_ _01679_ _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07944__A2 net483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09712_ _00291_ clknet_leaf_102_sys_clock_i internal_ih.received_byte_count\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07973_ net498 _03542_ _03543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06924_ _02442_ _02558_ _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA_hold464_I ci_neuron.uut_simple_neuron.titan_id_5\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08829__S _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09536__I3 _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06855_ _02081_ _02490_ _02491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09643_ ci_neuron.stream_o\[23\] net320 _04816_ _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05806_ _01058_ _01384_ _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09574_ _04768_ _04778_ _04779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06786_ _02372_ _02398_ _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold729_I _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08525_ _03785_ _04006_ _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05737_ _01304_ _01355_ _01401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06132__A1 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05668_ _01185_ _01187_ _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05052__I _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08456_ _01848_ _03948_ _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07407_ _02436_ _02454_ _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08387_ _03875_ _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07338_ _01946_ _01989_ _01991_ _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_05599_ ci_neuron.uut_simple_neuron.x2\[18\] _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_8_0_sys_clock_i clknet_0_sys_clock_i clknet_4_8_0_sys_clock_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_33_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07269_ _02898_ _01848_ _02713_ _02313_ _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_115_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09008_ _04355_ _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10280_ _00573_ clknet_leaf_129_sys_clock_i ci_neuron.stream_o\[22\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06199__B2 _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08538__I _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_81_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09369__I _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08974__I1 internal_ih.byte6\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_04970_ _00678_ _00034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_139_Right_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06640_ _02232_ _02280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_91_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06571_ _02210_ _02211_ _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05522_ ci_neuron.uut_simple_neuron.x2\[15\] ci_neuron.uut_simple_neuron.x2\[16\]
+ ci_neuron.uut_simple_neuron.x2\[17\] _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__09300__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09290_ net60 _04549_ _04555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08310_ _03825_ _03821_ _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05453_ _01117_ _01120_ _01122_ _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_08241_ _03761_ _03764_ _03765_ _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05384_ _00940_ _01055_ _01056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08172_ net680 net791 _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07123_ _02217_ _02237_ _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07614__A1 ci_neuron.uut_simple_neuron.x3\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07054_ _02678_ _02684_ _02686_ _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_88_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06005_ _01616_ _01663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_hold679_I _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08590__A2 _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07956_ _03512_ _03513_ _03527_ _03528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_126_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06907_ _02222_ _02506_ _02541_ _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_52_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07887_ _03457_ _03458_ _03470_ _03471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06838_ _02431_ _02458_ _02473_ _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09626_ _03926_ _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06769_ _02351_ _02353_ _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_108_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09557_ _04743_ _04759_ _04763_ _04764_ _00543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_93_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08508_ _03950_ _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09488_ _04697_ _04699_ _04703_ _04706_ _00532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_136_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08439_ _03939_ _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_137_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08653__I0 _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07081__A2 _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10263_ _00556_ clknet_leaf_98_sys_clock_i ci_neuron.stream_o\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10194_ _00120_ clknet_leaf_60_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05083__A1 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08947__I1 internal_ih.byte5\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07810_ ci_neuron.uut_simple_neuron.titan_id_4\[28\] ci_neuron.uut_simple_neuron.titan_id_3\[28\]
+ ci_neuron.uut_simple_neuron.titan_id_4\[27\] ci_neuron.uut_simple_neuron.titan_id_3\[27\]
+ _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08790_ _04027_ _01006_ _04225_ _04230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07741_ net582 _00103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04953_ internal_ih.byte0\[3\] _00665_ _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07672_ _03290_ _03291_ _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04884_ _00626_ _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06623_ _01883_ _02217_ _02263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09411_ _03754_ net60 _00814_ _01959_ _04622_ _04623_ _04640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_121_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06554_ _02180_ _02195_ _02196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_90_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09342_ _04584_ _00508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout30_I net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05505_ _01042_ _01173_ _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09890__CLK net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06485_ _02127_ _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09273_ _04543_ _04544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09380__S0 _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05436_ _01059_ _01106_ _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08224_ _03747_ _03750_ _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_117_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05367_ _00976_ _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08155_ net684 ci_neuron.uut_simple_neuron.titan_id_0\[26\] _03693_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07106_ _02737_ _02617_ _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_76_sys_clock_i clknet_4_10_0_sys_clock_i clknet_leaf_76_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05298_ _00971_ _00964_ _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08086_ net519 _03636_ _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07037_ _02614_ _02630_ _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09472__I _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08988_ _04343_ _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07939_ _03512_ net571 _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_3_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05129__A2 _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09609_ net351 ci_neuron.output_memory\[8\] _04800_ _04801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04888__A1 internal_ih.byte4\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06629__A2 _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09418__I2 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10246_ _00143_ clknet_leaf_17_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10177_ _00074_ clknet_leaf_119_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06270_ _01909_ _01911_ _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08490__A1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_96_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05221_ _00894_ _00897_ _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xclkbuf_leaf_118_sys_clock_i clknet_4_6_0_sys_clock_i clknet_leaf_118_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_7_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold615 ci_neuron.uut_simple_neuron.titan_id_3\[26\] net648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold604 ci_neuron.uut_simple_neuron.titan_id_3\[14\] net637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05152_ _00784_ _00821_ _00823_ _00810_ _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
Xhold626 ci_neuron.uut_simple_neuron.titan_id_5\[16\] net659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_69_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05083_ _00749_ _00754_ _00764_ _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold637 ci_neuron.uut_simple_neuron.titan_id_0\[18\] net670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold659 _03677_ net692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold648 _03705_ net681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09960_ _00475_ clknet_leaf_3_sys_clock_i ci_neuron.uut_simple_neuron.x0\[31\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08911_ net496 _00362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09891_ _00052_ net18 ci_neuron.value_i\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold377_I internal_ih.byte4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08842_ _04170_ _04254_ _04260_ _00332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_99_sys_clock_i_I clknet_4_10_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05985_ _01492_ _01547_ _01548_ _01641_ _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08773_ _00814_ _04214_ _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07724_ _03334_ net638 _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_0_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04936_ _00626_ _00659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07655_ net713 ci_neuron.uut_simple_neuron.titan_id_3\[2\] _03278_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06606_ _02204_ _02203_ _02247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_105_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04867_ internal_ih.byte7\[3\] _00606_ _00614_ _00610_ _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07586_ _03152_ _03211_ _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06537_ _02178_ _02146_ _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09325_ _04074_ net75 _04572_ _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06468_ _02073_ _02108_ _02111_ _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_90_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_25_sys_clock_i clknet_4_6_0_sys_clock_i clknet_leaf_25_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09256_ _04122_ net551 _04490_ _04532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05419_ _01018_ _01046_ _01089_ _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_60_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08207_ net170 net163 _03736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_134_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06399_ _02000_ _02044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_62_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09187_ _00706_ _04491_ _04493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08138_ net691 ci_neuron.uut_simple_neuron.titan_id_0\[22\] _03679_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08069_ _03618_ _03619_ _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_116_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10100_ _00166_ clknet_leaf_55_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05598__A2 _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10031_ net181 clknet_leaf_94_sys_clock_i ci_neuron.output_val_internal\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05286__B2 _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10229_ _00156_ clknet_leaf_87_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05770_ net760 _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07440_ _02993_ _03055_ _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07371_ _02926_ _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06322_ _01968_ _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_128_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09110_ net139 _04416_ _04450_ _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_33_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08463__A1 _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09041_ _04383_ ci_neuron.stream_o\[1\] ci_neuron.stream_o\[17\] _04384_ _04387_
+ _04388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_111_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06253_ _01872_ _01879_ _01901_ _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_103_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09287__I _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_87_sys_clock_i_I clknet_4_11_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06184_ _01835_ _01836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05204_ _00818_ _00880_ _00872_ _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08215__A1 _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold401 internal_ih.byte7\[2\] net434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold412 ci_neuron.uut_simple_neuron.titan_id_4\[24\] net445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_130_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold423 ci_neuron.uut_simple_neuron.titan_id_4\[13\] net456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05135_ _00753_ _00793_ _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold445 internal_ih.byte0\[7\] net478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold434 _04297_ net467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_hold494_I internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold467 ci_neuron.input_memory\[1\]\[6\] net628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold478 ci_neuron.uut_simple_neuron.x0\[5\] net511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold456 internal_ih.byte2\[7\] net489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_110_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold489 _03300_ net522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05066_ _00749_ _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09943_ _00458_ clknet_leaf_117_sys_clock_i ci_neuron.uut_simple_neuron.x0\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_hold661_I _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09874_ _00034_ net28 ci_neuron.value_i\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08825_ _04110_ _01792_ _04246_ _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_135_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05968_ _01526_ _01626_ _01627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05055__I _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08756_ _04208_ _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_49_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05899_ _01557_ _01541_ _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07707_ _03312_ _03318_ _03321_ _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08687_ _04134_ _04151_ _04153_ _00284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04919_ internal_ih.byte5\[5\] _00646_ _00647_ internal_ih.byte1\[5\] _00649_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_138_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07638_ _03261_ _03262_ _03263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07569_ _03126_ _03128_ _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08829__I0 _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09308_ _04034_ net80 _04561_ _04565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08454__A1 ci_neuron.value_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09239_ _04085_ _03864_ _04519_ _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_134_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09254__I0 _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_79_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_73_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10014_ net80 clknet_leaf_48_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08693__B2 _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10193__D _00118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_97_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06940_ _02519_ _02518_ _02574_ _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06871_ _02222_ _02506_ _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input2_I spi_cs_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05822_ _01428_ _01429_ _01483_ _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08610_ _04087_ _00273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09590_ _04789_ _04790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05753_ _01369_ _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08541_ _04027_ _02228_ _04028_ _04029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05684_ _01323_ _01348_ _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_82_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08472_ _03967_ _01872_ _03969_ _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07423_ _01892_ _03050_ _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08684__B2 _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09079__I3 ci_neuron.output_val_internal\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07354_ _02981_ _02843_ _02982_ _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_118_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07239__A2 ci_neuron.uut_simple_neuron.x3\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08914__I _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout7_I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07285_ _02845_ _02914_ _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06305_ _01829_ _01876_ _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06236_ _01836_ _01839_ _01865_ _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09024_ net206 _04354_ _04371_ _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_131_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold220 net4 net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_06167_ ci_neuron.uut_simple_neuron.x3\[1\] _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold242 _01266_ net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold231 ci_neuron.uut_simple_neuron.titan_id_6\[8\] net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold253 internal_ih.current_instruction\[4\] net286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_113_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold264 _03294_ net297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05118_ _00790_ _00798_ _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold286 _01754_ net319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_06098_ ci_neuron.uut_simple_neuron.x2\[27\] _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold275 _04797_ net308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05049_ _00733_ _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold297 _03887_ net330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09926_ _00031_ net5 ci_neuron.instruction_i\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_129_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07175__A1 _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_144_sys_clock_i_I clknet_4_0_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09857_ _00436_ clknet_leaf_125_sys_clock_i ci_neuron.output_memory\[25\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08808_ _04069_ net550 _04239_ _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09788_ _00367_ clknet_leaf_142_sys_clock_i internal_ih.byte4\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_142_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08739_ _04193_ _04196_ _04197_ _00292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_142_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08427__A1 _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09490__I3 _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_75_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09390__I _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08734__I _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07070_ _02644_ _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06021_ _01654_ _01678_ _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_63_sys_clock_i_I clknet_4_15_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09394__A2 _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold192_I ci_neuron.output_val_internal\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09711_ net185 clknet_leaf_105_sys_clock_i spi_interface_cvonk.buffer\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07972_ net786 net624 _03542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06923_ _02554_ _02557_ _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_06854_ _02053_ _02489_ _02490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09642_ net299 _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06785_ _02419_ _02421_ _02422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05805_ _01208_ _01389_ _01466_ _01467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09573_ _03916_ ci_neuron.input_memory\[1\]\[30\] _01793_ ci_neuron.uut_simple_neuron.x3\[30\]
+ _04760_ _04761_ _04778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_132_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05736_ _01396_ _01399_ _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08524_ _04005_ _03998_ _03783_ _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_78_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05667_ _01186_ _01287_ _01223_ _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08455_ _00065_ _03952_ _03954_ _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07406_ _03032_ _03033_ _03034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05598_ _01227_ _01264_ _01265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07880__A2 ci_neuron.uut_simple_neuron.titan_id_5\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08386_ _03891_ _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07337_ _02964_ _02965_ _02966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_132_sys_clock_i_I clknet_4_2_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07268_ _01847_ _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_103_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07199_ _02827_ _02829_ _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06219_ _01858_ _01868_ _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09007_ _04177_ _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09909_ _00005_ net9 ci_neuron.address_i\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05634__A1 _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06570_ _01889_ _02176_ _02211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_51_sys_clock_i_I clknet_4_13_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05521_ _01097_ _01149_ _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_87_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09300__A2 _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05452_ _01074_ _01077_ _01115_ _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_90_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ net596 net763 _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_145_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05873__A1 _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08171_ _03706_ _00084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07122_ _02752_ _02753_ _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_99_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05383_ _01053_ _01054_ _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07614__A2 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07053_ _02379_ _02685_ _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05625__A1 _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06004_ _01617_ _01623_ _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06050__A1 _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07955_ ci_neuron.uut_simple_neuron.titan_id_2\[19\] ci_neuron.uut_simple_neuron.titan_id_5\[19\]
+ _03527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_52_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_126_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06906_ _02223_ _02379_ _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_52_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07145__A4 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07886_ _03453_ _03460_ _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09625_ net365 _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06837_ _02434_ _02457_ _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06353__A2 _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_120_sys_clock_i_I clknet_4_3_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06768_ _02405_ _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_108_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09556_ net186 _04749_ _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06699_ ci_neuron.uut_simple_neuron.x3\[15\] ci_neuron.uut_simple_neuron.x3\[16\]
+ _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05719_ _01344_ _01328_ _01382_ _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08507_ _03770_ _03987_ _03772_ _03999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09487_ net144 _04705_ _04706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08438_ _03938_ _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_43_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08369_ _03874_ _03877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10262_ _00555_ clknet_leaf_98_sys_clock_i ci_neuron.stream_o\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_52_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10193_ _00118_ clknet_leaf_91_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06041__A1 _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06344__A2 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07541__A1 _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09294__A1 _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_117_sys_clock_i clknet_4_9_0_sys_clock_i clknet_leaf_117_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_25_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07740_ _03347_ _03348_ _03349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04952_ _00668_ _00055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07671_ _03287_ _03288_ _03291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04883_ _00603_ _00596_ _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06622_ _02213_ _02260_ _02261_ _02262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09410_ ci_neuron.output_memory\[6\] _04628_ _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_121_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06553_ _02194_ _02191_ _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09341_ _04110_ net93 _04583_ _04584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05504_ _00981_ _01140_ _01173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06484_ _01896_ _01994_ _02126_ _02127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_24_sys_clock_i clknet_4_6_0_sys_clock_i clknet_leaf_24_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09272_ _04542_ _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09380__S1 _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05435_ _01098_ _01105_ _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08223_ _03748_ _03749_ _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05366_ _00972_ _01035_ _01037_ _01038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08154_ _03688_ net743 _03691_ _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__09588__A2 _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07599__A1 _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07105_ _02736_ _02733_ _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08085_ _03635_ _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07036_ _02614_ _02630_ _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05297_ _00970_ _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05058__I _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08987_ _04146_ _00594_ _04339_ _04343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07938_ ci_neuron.uut_simple_neuron.titan_id_2\[19\] net570 _03513_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07869_ _03429_ _03432_ _03454_ _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09608_ _04789_ _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09539_ net233 _04749_ _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09418__I3 _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09579__A2 _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_60_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09200__A1 _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10245_ _00142_ clknet_leaf_17_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10176_ _00073_ clknet_leaf_119_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08279__I _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09503__A2 _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08562__I0 _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05220_ _00740_ _00896_ _00897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_96_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05151_ _00806_ _00827_ _00829_ _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold616 _03396_ net649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold605 _03335_ net638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold627 _03504_ net660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_123_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06253__A1 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05082_ _00733_ _00753_ _00757_ _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xhold649 ci_neuron.input_memory\[1\]\[20\] net757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold638 _03664_ net671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_1_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08910_ internal_ih.byte4\[0\] net495 _04296_ _04299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09890_ _00051_ net23 ci_neuron.value_i\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08841_ internal_ih.byte0\[2\] _04254_ _04260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_85_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05984_ _01550_ _01641_ _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08772_ _03979_ _04218_ _04219_ _00303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07505__A1 _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_108_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07723_ ci_neuron.uut_simple_neuron.titan_id_4\[14\] net637 _03335_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_0_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04935_ _00639_ _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_hold537_I ci_neuron.uut_simple_neuron.titan_id_5\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07654_ net713 ci_neuron.uut_simple_neuron.titan_id_3\[2\] _03277_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_0_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06605_ _02245_ _02202_ _02246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04866_ internal_ih.byte4\[3\] internal_ih.byte3\[3\] _00608_ _00614_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07585_ _03155_ _03210_ _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06536_ _02138_ _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09324_ _04574_ _00500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06467_ _01985_ _02109_ _02110_ _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_118_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09255_ _04531_ _00474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Left_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05418_ _00940_ _01011_ _01007_ _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08206_ net32 net170 net163 _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06398_ _02006_ _02010_ _02042_ _02043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_90_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09186_ _03947_ _04489_ _04492_ _00444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_134_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07268__I _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05349_ _01010_ _01021_ _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08137_ ci_neuron.uut_simple_neuron.titan_id_1\[22\] ci_neuron.uut_simple_neuron.titan_id_0\[22\]
+ _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_141_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06244__A1 _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06172__I ci_neuron.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08068_ ci_neuron.uut_simple_neuron.titan_id_1\[10\] ci_neuron.uut_simple_neuron.titan_id_0\[10\]
+ _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07019_ _02593_ _02650_ _02651_ _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_116_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10030_ _00515_ clknet_leaf_110_sys_clock_i internal_ih.data_pointer\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_126_Left_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_135_Left_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_144_Left_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08511__B _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10228_ _00155_ clknet_leaf_87_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10159_ net65 clknet_leaf_92_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08535__I0 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08160__A1 _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07370_ _02950_ _02960_ _02997_ _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06321_ _01967_ _01896_ _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_45_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06252_ _01873_ _01900_ _01901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_100_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09040_ _04385_ _04386_ _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05203_ _00751_ _00842_ _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06183_ _01834_ _01835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold402 _04333_ net435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_142_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold413 _03387_ net446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_111_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06226__A1 _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold424 _03331_ net457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05134_ _00813_ _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold435 internal_ih.byte1\[1\] net468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_05065_ _00748_ _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09942_ _00457_ clknet_leaf_71_sys_clock_i ci_neuron.uut_simple_neuron.x0\[13\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold468 internal_ih.byte0\[1\] net501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold446 _04277_ net479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold457 _04298_ net490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold479 _03751_ net512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06720__I _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09873_ _00064_ net27 ci_neuron.value_i\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08824_ net319 _04236_ _04249_ _00325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08755_ _04207_ _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05967_ _01611_ _01625_ _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07706_ _03319_ _03320_ _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05898_ _01557_ _01541_ _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08686_ _04152_ _04149_ _04153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04918_ _00648_ _00004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__04960__A1 internal_ih.byte0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07637_ _03197_ _03208_ _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04849_ _00594_ _00599_ _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07568_ _03157_ _03193_ _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_62_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06519_ _02158_ _02161_ _02162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09307_ _04564_ _00493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07499_ _03124_ _03125_ _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09478__I _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08454__A2 _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09238_ _04079_ _04503_ _04522_ _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_51_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09169_ net232 _04481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09254__I1 _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10013_ net74 clknet_leaf_71_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04951__A1 internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ _02188_ _02337_ _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05821_ _01368_ _01381_ _01480_ _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_89_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05752_ _01412_ _01391_ _01414_ _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08540_ _03968_ _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_77_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05683_ _01218_ _01325_ _01347_ _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_08471_ _03968_ _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07422_ _03047_ _03049_ _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07353_ _02913_ _02982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_118_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07284_ _02846_ _02913_ _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06304_ _01949_ _01937_ _01950_ _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_118_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06235_ _01827_ _01884_ _01885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_60_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09023_ _04356_ _04364_ _04369_ _04370_ _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_131_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold210 ci_neuron.uut_simple_neuron.titan_id_6\[20\] net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06166_ _01819_ _01820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold232 ci_neuron.uut_simple_neuron.titan_id_6\[14\] net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold221 _04132_ net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold243 ci_neuron.output_memory\[17\] net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_113_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05117_ _00734_ _00792_ _00797_ _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_06097_ _01750_ _01752_ _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_hold771_I internal_ih.byte1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold276 ci_neuron.output_memory\[4\] net309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold265 ci_neuron.output_memory\[22\] net298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold287 ci_neuron.output_memory\[23\] net320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold254 ci_neuron.uut_simple_neuron.titan_id_0\[2\] net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_102_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05048_ net33 _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold298 _03888_ net331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09925_ _00030_ net11 ci_neuron.instruction_i\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09856_ _00435_ clknet_leaf_124_sys_clock_i ci_neuron.output_memory\[24\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07175__A2 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05066__I _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08807_ _04240_ _00317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06999_ _02606_ _02632_ _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_99_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09787_ _00366_ clknet_leaf_141_sys_clock_i internal_ih.byte4\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_142_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08738_ net293 _04195_ _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08669_ _04136_ _04137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06686__A1 _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08427__A2 _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09001__I net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07456__I _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06677__A1 _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08910__I0 internal_ih.byte4\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_74_sys_clock_i clknet_4_12_0_sys_clock_i clknet_leaf_74_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06020_ _01568_ _01677_ _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07971_ net825 net497 _03530_ _03538_ _03540_ _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06922_ _02498_ _02556_ _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09710_ net132 clknet_leaf_105_sys_clock_i internal_ih.spi_rx_byte_i\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06853_ _02181_ _02453_ _02488_ _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_93_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09641_ ci_neuron.stream_o\[22\] net298 _04816_ _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06784_ _02420_ _02368_ _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05804_ _01462_ _01463_ _01465_ _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09572_ ci_neuron.output_memory\[30\] _04766_ _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05735_ _01397_ _01398_ _01399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08523_ _04000_ _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08901__I0 internal_ih.byte3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05666_ _01292_ _01293_ _01330_ _01268_ _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_08454_ ci_neuron.value_i\[1\] _03953_ _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07969__C net458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07405_ _02382_ _02947_ _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05597_ ci_neuron.uut_simple_neuron.x2\[19\] _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08385_ ci_neuron.uut_simple_neuron.x0\[27\] _03891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07336_ _02888_ _02894_ _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07267_ _02852_ _02896_ _02897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_131_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09006_ _04182_ _04354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07198_ _01907_ _02828_ _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_131_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06840__A1 _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06218_ _01860_ _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06149_ _01743_ _01796_ _01803_ _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_57_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09908_ _00004_ net9 ci_neuron.address_i\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09839_ _00418_ clknet_leaf_89_sys_clock_i ci_neuron.output_memory\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05331__A1 _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_116_sys_clock_i clknet_4_9_0_sys_clock_i clknet_leaf_116_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09620__I1 ci_neuron.output_memory\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05570__A1 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05520_ _01147_ _01151_ _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_23_sys_clock_i clknet_4_6_0_sys_clock_i clknet_leaf_23_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05451_ _01121_ _00206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08170_ _03704_ net681 _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07075__A1 _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07121_ _02184_ _02691_ _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05382_ ci_neuron.uut_simple_neuron.x2\[12\] ci_neuron.uut_simple_neuron.x2\[13\]
+ ci_neuron.uut_simple_neuron.x2\[14\] _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_15_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07052_ _02339_ _02500_ _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_88_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06003_ _01462_ _01660_ _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09611__I1 ci_neuron.output_memory\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06050__A2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07954_ _03518_ _03523_ _03526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06905_ _02491_ _02510_ _02539_ _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_126_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07885_ _03462_ _03465_ _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06836_ _02470_ _02471_ _02472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09624_ net364 ci_neuron.output_memory\[15\] _04805_ _04809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06767_ _02401_ _02404_ _02405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_108_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09555_ _04746_ _04762_ _04763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06698_ _02228_ _02334_ _02336_ _02337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05718_ _01342_ _01381_ _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08506_ _03997_ _03998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09486_ _04704_ _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05649_ _01304_ _01314_ _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_109_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08437_ _03933_ _03937_ _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08368_ _03874_ _03875_ _03876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07319_ _02382_ _02947_ _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08299_ _03804_ _03805_ _03815_ _03803_ _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_103_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09486__I _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10261_ _00554_ clknet_leaf_98_sys_clock_i ci_neuron.stream_o\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08566__A1 _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10192_ _00107_ clknet_leaf_91_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08766__S _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05552__A1 _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09396__I _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08557__A1 _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04951_ internal_ih.byte0\[2\] _00665_ _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07670_ ci_neuron.uut_simple_neuron.titan_id_4\[5\] ci_neuron.uut_simple_neuron.titan_id_3\[5\]
+ _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04882_ _00605_ _00625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06621_ _02215_ _02240_ _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05543__A1 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06552_ _02193_ _02194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_87_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09340_ _04566_ _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05503_ _01144_ _01154_ _01171_ _01132_ _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_90_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09285__A2 _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09271_ _03933_ _04485_ _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_47_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06483_ _02100_ _02101_ _02126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08222_ _03729_ net511 net173 _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_05434_ _01104_ _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05365_ _01036_ _01021_ _01037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08153_ net742 net792 _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07104_ _02735_ _02734_ _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08084_ ci_neuron.uut_simple_neuron.titan_id_1\[13\] ci_neuron.uut_simple_neuron.titan_id_0\[13\]
+ _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07035_ _02661_ _02667_ _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05296_ _00969_ _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_54_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08986_ _00598_ _04340_ _04342_ _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07937_ _03508_ _03509_ _03511_ _03512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_138_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07868_ ci_neuron.uut_simple_neuron.titan_id_2\[3\] ci_neuron.uut_simple_neuron.titan_id_5\[3\]
+ _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06819_ _02452_ _02455_ _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07799_ net649 net783 _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09607_ net312 _00558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09538_ _04704_ _04749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09276__A2 _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09469_ _04673_ _04686_ _04688_ _04689_ _00530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_93_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10244_ _00141_ clknet_leaf_124_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07211__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10175_ _00072_ clknet_leaf_23_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08562__I1 _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07278__A1 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05150_ _00802_ _00825_ _00824_ _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08778__A1 _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold606 _03336_ net639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_69_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold617 ci_neuron.input_memory\[1\]\[27\] net714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_122_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05081_ _00735_ _00761_ _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold639 ci_neuron.uut_simple_neuron.titan_id_1\[11\] net672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold628 ci_neuron.uut_simple_neuron.titan_id_2\[2\] net661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09578__I0 ci_neuron.uut_simple_neuron.x0\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08840_ _04259_ _00331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05983_ _01597_ _01637_ _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_109_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08771_ net829 _04214_ _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07722_ _03330_ _03332_ _03333_ _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_0_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04934_ _00657_ _00011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07653_ net653 _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04865_ _00613_ _00027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06604_ _02199_ _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_105_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07584_ _03194_ _03209_ _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_125_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09323_ _04069_ net77 _04572_ _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07269__A1 _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06535_ _01856_ _02176_ _02177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06466_ _02036_ _02061_ _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ _04119_ _03916_ _04490_ _04531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_106_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05417_ _01083_ _01086_ _01087_ _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08205_ _03729_ _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09185_ _03725_ _04491_ _04492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06397_ _02040_ _02041_ _02042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08769__A1 _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08136_ net692 _00078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05348_ _01012_ _01000_ _01020_ _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__06244__A2 _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05279_ _00952_ _00953_ _00954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_70_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08067_ net726 _00094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07018_ _02596_ _02633_ _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_116_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09682__CLK clknet_4_7_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08969_ _04192_ _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_27_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09004__I _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10227_ _00154_ clknet_leaf_90_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10158_ net66 clknet_leaf_78_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10089_ _00186_ clknet_leaf_10_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[26\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08535__I1 _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06320_ _01963_ net164 _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_85_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06251_ _01878_ _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_100_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05202_ _00855_ _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_53_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06182_ ci_neuron.uut_simple_neuron.x3\[0\] _01822_ _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09412__A2 _04640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07423__A1 _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05133_ _00812_ _00813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold425 ci_neuron.uut_simple_neuron.titan_id_5\[22\] net458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold414 ci_neuron.input_memory\[1\]\[5\] net597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold403 ci_neuron.uut_simple_neuron.x0\[28\] net436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold436 _04279_ net469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05064_ _00747_ _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xhold447 ci_neuron.uut_simple_neuron.x2\[31\] net480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09941_ _00456_ clknet_leaf_116_sys_clock_i ci_neuron.uut_simple_neuron.x0\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold458 internal_ih.byte4\[1\] net491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold469 net813 net502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09872_ _00063_ net29 ci_neuron.value_i\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08823_ _04104_ _04237_ _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05966_ _01616_ _01624_ _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08754_ _03937_ _04206_ _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07705_ ci_neuron.uut_simple_neuron.titan_id_4\[10\] ci_neuron.uut_simple_neuron.titan_id_3\[10\]
+ net411 net598 _03320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_04917_ internal_ih.byte5\[4\] _00646_ _00647_ internal_ih.byte1\[4\] _00648_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05897_ _01252_ _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_49_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08685_ internal_ih.spi_rx_byte_i\[2\] _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07636_ _03200_ _03207_ _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04848_ _00598_ internal_ih.current_instruction\[3\] internal_ih.current_instruction\[2\]
+ _00592_ _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_138_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07567_ _03181_ _03192_ _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06518_ _02073_ _02159_ _02160_ _02161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09306_ _04027_ net74 _04561_ _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07498_ _01984_ _03048_ _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09237_ _03862_ _04496_ _04522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06449_ _01998_ _02050_ _02092_ _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_106_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_59_sys_clock_i_I clknet_4_14_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09168_ _04480_ _00438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08119_ _03662_ _03663_ _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09099_ _04365_ _04440_ _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07965__A2 ci_neuron.uut_simple_neuron.titan_id_5\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10012_ net96 clknet_leaf_70_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08838__I _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05262__I _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_73_sys_clock_i clknet_4_9_0_sys_clock_i clknet_leaf_73_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_54_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_128_sys_clock_i_I clknet_4_3_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07405__A1 _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05820_ _01477_ _01481_ _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05751_ _01413_ _01390_ _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05682_ _01331_ _01341_ _01346_ _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08470_ _03938_ _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07421_ _01984_ _03048_ _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_106_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07352_ _02846_ _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_119_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06303_ _01928_ _01948_ _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07283_ _02910_ _02912_ _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_115_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06234_ _01871_ _01883_ _01884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_60_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09022_ _04182_ _04370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_131_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06165_ ci_neuron.uut_simple_neuron.x3\[0\] _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold200 ci_neuron.output_val_internal\[24\] net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold211 ci_neuron.output_val_internal\[31\] net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05116_ _00794_ _00796_ _00797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07947__A2 net483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold222 _00282_ net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_14_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold244 _04813_ net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold233 ci_neuron.uut_simple_neuron.titan_id_6\[1\] net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_141_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06096_ _00937_ _01751_ _01669_ _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold277 _04796_ net310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold266 _04819_ net299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold255 _03723_ net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09924_ _00029_ net5 ci_neuron.instruction_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold288 _04820_ net321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold299 ci_neuron.stream_o\[14\] net332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05047_ _00715_ _00725_ _00732_ _00000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09855_ _00434_ clknet_leaf_120_sys_clock_i ci_neuron.output_memory\[23\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08806_ _04064_ net762 _04239_ _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06998_ _02631_ _02608_ _02632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09786_ _00365_ clknet_leaf_137_sys_clock_i internal_ih.byte4\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_134_Right_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05949_ _01576_ _01585_ _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_47_sys_clock_i_I clknet_4_6_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08737_ net293 _04195_ _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_139_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08668_ _04135_ _04136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_37_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07619_ _03181_ _03192_ _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08599_ _04076_ _04077_ _03953_ _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_49_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_115_sys_clock_i clknet_4_9_0_sys_clock_i clknet_leaf_115_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_106_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07938__A2 net570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05257__I _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_116_sys_clock_i_I clknet_4_9_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09560__A1 net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_86_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_22_sys_clock_i clknet_4_6_0_sys_clock_i clknet_leaf_22_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09399__I _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07970_ _03539_ _03540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06921_ ci_neuron.uut_simple_neuron.x3\[19\] _02555_ _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__09551__A1 ci_neuron.output_memory\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06852_ _02182_ _02329_ _02488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09640_ net472 _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06783_ _01920_ _01938_ _02420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05803_ _01464_ _01431_ _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09571_ _04765_ _04773_ _04775_ _04776_ _00545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05734_ _00932_ _01351_ _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08522_ _03986_ _04010_ _04012_ _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08453_ _03925_ _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09893__CLK net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07404_ _02392_ _02946_ _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05665_ _00936_ _01329_ _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_46_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05596_ _01099_ _01102_ _01187_ _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_73_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08384_ _03889_ _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07335_ _02891_ _02893_ _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07266_ _02885_ _02895_ _02896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06217_ _01823_ _01867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09005_ _04351_ _04353_ _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07197_ _02273_ _02291_ _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_35_sys_clock_i_I clknet_4_5_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06148_ _01621_ _01802_ _01803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_57_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06079_ _01648_ _01725_ _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08593__A2 _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09907_ _00003_ net10 ci_neuron.address_i\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09838_ _00417_ clknet_leaf_88_sys_clock_i ci_neuron.output_memory\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09769_ _00348_ clknet_leaf_138_sys_clock_i internal_ih.byte2\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06108__A1 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09012__I internal_ih.data_pointer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07084__A2 _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_104_sys_clock_i_I clknet_4_8_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05450_ _01118_ _01120_ _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05381_ _00970_ _01005_ _01052_ _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08647__I0 _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07120_ _02190_ _02690_ _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_99_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07051_ _02502_ _02683_ _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_70_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06281__I _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06002_ _01374_ _01659_ _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_51_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold295_I ci_neuron.output_memory\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07953_ ci_neuron.uut_simple_neuron.titan_id_2\[21\] net414 _03525_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06904_ _02493_ _02509_ _02539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07884_ ci_neuron.uut_simple_neuron.titan_id_2\[9\] ci_neuron.uut_simple_neuron.titan_id_5\[9\]
+ _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_52_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold462_I internal_ih.byte3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06835_ _02365_ _02430_ _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09623_ net333 _00565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06766_ _02266_ _02402_ _02403_ _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_108_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09554_ _03892_ ci_neuron.input_memory\[1\]\[27\] _01706_ _03084_ _04760_ _04761_
+ _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_06697_ _02335_ _02333_ _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05717_ net738 _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_23_sys_clock_i_I clknet_4_6_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08505_ _03769_ _03771_ _03987_ _03997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09485_ _04596_ _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05648_ _01313_ _01314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08436_ _03934_ _03936_ _03937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08367_ net329 _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07318_ _02392_ _02946_ _02947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05579_ _01246_ _00209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08298_ net347 ci_neuron.uut_simple_neuron.x0\[15\] _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07249_ _02878_ _02857_ _02879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_10260_ _00553_ clknet_leaf_98_sys_clock_i ci_neuron.stream_o\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06577__A1 _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08810__I0 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10191_ _00096_ clknet_leaf_92_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08782__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09054__I0 ci_neuron.output_val_internal\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04950_ _00667_ _00044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06620_ _02215_ _02240_ _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_04881_ _00624_ _00032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_87_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08756__I _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06551_ _01954_ _02192_ _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06482_ _01846_ _02125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05502_ _01058_ _01152_ _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09270_ _04540_ _04535_ net301 _00479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05433_ _01103_ _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08221_ net173 net511 _03733_ _03737_ _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_8_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07048__A2 ci_neuron.uut_simple_neuron.x3\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05364_ _01010_ _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08152_ _03690_ _00081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_136_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07103_ _02730_ ci_neuron.uut_simple_neuron.x3\[23\] _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_05295_ ci_neuron.uut_simple_neuron.x2\[12\] _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08083_ net518 ci_neuron.uut_simple_neuron.titan_id_0\[12\] _03631_ _03632_ _03634_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07034_ _02664_ _02666_ _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09045__I0 ci_neuron.output_val_internal\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06559__A1 _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_11_sys_clock_i_I clknet_4_4_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08985_ _04143_ _04341_ _04342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07936_ ci_neuron.uut_simple_neuron.titan_id_2\[18\] ci_neuron.uut_simple_neuron.titan_id_5\[18\]
+ _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07867_ ci_neuron.uut_simple_neuron.titan_id_2\[7\] ci_neuron.uut_simple_neuron.titan_id_5\[7\]
+ _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06818_ _02454_ _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07798_ net782 ci_neuron.uut_simple_neuron.titan_id_3\[27\] _03397_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09606_ ci_neuron.stream_o\[7\] net311 _04795_ _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06749_ ci_neuron.uut_simple_neuron.x3\[15\] _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09537_ _04746_ _04747_ _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_65_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_6_sys_clock_i_I clknet_4_4_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09468_ net115 _04680_ _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_22_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09399_ _04602_ _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08419_ _03919_ _03920_ _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_123_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10243_ _00140_ clknet_leaf_120_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10174_ _00071_ clknet_leaf_70_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold607 ci_neuron.uut_simple_neuron.titan_id_4\[22\] net640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold618 ci_neuron.uut_simple_neuron.x0\[21\] net744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_05080_ _00758_ _00759_ _00762_ _00161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold629 _03426_ net662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_122_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05213__A1 _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05982_ _01640_ _00218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08770_ _04208_ _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_9_sys_clock_i clknet_4_4_0_sys_clock_i clknet_leaf_9_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07721_ net456 ci_neuron.uut_simple_neuron.titan_id_3\[13\] _03333_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04933_ internal_ih.byte6\[3\] _00652_ _00653_ internal_ih.byte2\[3\] _00657_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07652_ ci_neuron.uut_simple_neuron.titan_id_4\[2\] ci_neuron.uut_simple_neuron.titan_id_3\[2\]
+ _03275_ _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_0_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04864_ internal_ih.byte7\[2\] _00606_ _00612_ _00610_ _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07583_ _03197_ _03208_ _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06603_ _02241_ _02243_ _02244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_105_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06534_ _01862_ _02175_ _02176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09322_ _04573_ _00499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07269__A2 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold425_I ci_neuron.uut_simple_neuron.titan_id_5\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08466__A1 _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06465_ _02036_ _02061_ _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09253_ _04530_ _00473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_145_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06396_ _02005_ _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_105_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05416_ _01084_ _01085_ _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_62_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08204_ net528 net173 _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09184_ _04490_ _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05347_ _01018_ _01019_ _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08135_ net691 ci_neuron.uut_simple_neuron.titan_id_0\[22\] _03676_ _03677_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_60_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05278_ _00931_ _00933_ _00950_ _00953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08066_ _03618_ net725 _03620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_141_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07017_ _02596_ _02633_ _02650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_116_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09194__A2 _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08968_ net340 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07919_ _03493_ _03495_ _03496_ _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_08899_ internal_ih.byte3\[3\] net269 _04291_ _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_27_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05507__A2 _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08457__A1 _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_72_sys_clock_i clknet_4_12_0_sys_clock_i clknet_leaf_72_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_35_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_49_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_132_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10226_ _00153_ clknet_leaf_90_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09185__A2 _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10157_ _00222_ clknet_leaf_35_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10088_ _00185_ clknet_leaf_11_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09488__A3 _04703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08448__A1 _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06250_ _01898_ _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09248__I0 _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05201_ _00851_ _00875_ _00877_ _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08970__S _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06181_ _01833_ _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05132_ _00811_ _00812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold415 ci_neuron.input_memory\[1\]\[9\] net626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold404 internal_ih.byte6\[0\] net437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold426 _03533_ net459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05063_ ci_neuron.uut_simple_neuron.x2\[1\] _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09940_ _00455_ clknet_leaf_116_sys_clock_i ci_neuron.uut_simple_neuron.x0\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold437 net814 net470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold448 net815 net481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold459 internal_ih.byte3\[7\] net492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_25_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09871_ _00062_ net29 ci_neuron.value_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08822_ _01619_ _04236_ _04248_ _00324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05965_ _01617_ _01623_ _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08753_ _03934_ _03931_ _03928_ _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07704_ ci_neuron.uut_simple_neuron.titan_id_4\[10\] ci_neuron.uut_simple_neuron.titan_id_3\[10\]
+ _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04916_ _00627_ _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05896_ _01518_ _01554_ _01555_ _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_49_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08684_ net161 _04137_ _04142_ _04146_ _04151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07635_ _03242_ _03245_ _03259_ _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_49_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04847_ net279 _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xclkbuf_leaf_114_sys_clock_i clknet_4_9_0_sys_clock_i clknet_leaf_114_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07566_ _03184_ _03191_ _03192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06517_ _02108_ _02111_ _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09305_ _04563_ _00492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07497_ _02040_ _02009_ _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09236_ _04521_ _00465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06448_ _02089_ _02091_ _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_106_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09239__I0 _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_32_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06379_ _01981_ _02024_ _02023_ _02025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09167_ net252 _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07414__A2 _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08118_ net663 ci_neuron.uut_simple_neuron.titan_id_0\[19\] _03663_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09098_ ci_neuron.output_val_internal\[30\] ci_neuron.output_val_internal\[22\] ci_neuron.output_val_internal\[14\]
+ ci_neuron.output_val_internal\[6\] _04366_ _04367_ _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08049_ net603 ci_neuron.uut_simple_neuron.titan_id_0\[7\] _03605_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07178__A1 _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10011_ net84 clknet_leaf_69_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06925__A1 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_21_sys_clock_i clknet_4_3_0_sys_clock_i clknet_leaf_21_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_57_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08790__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08602__A1 _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07169__A1 ci_neuron.uut_simple_neuron.x3\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10209_ _00105_ clknet_leaf_44_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_66_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05750_ _01208_ _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05681_ _01330_ _01343_ _01345_ _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_82_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07420_ _01997_ _02008_ _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07351_ _02840_ _02914_ _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_75_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06302_ _01928_ _01948_ _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_128_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07282_ _02781_ _02834_ _02911_ _02912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08841__A1 internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06233_ _01882_ _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09021_ _04365_ _04368_ _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_131_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06164_ _01818_ _00222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold201 _00540_ net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05115_ _00756_ _00766_ _00795_ _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xhold234 internal_ih.received_byte_count\[7\] net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold223 internal_ih.received_byte_count\[1\] net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09641__I0 ci_neuron.stream_o\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold212 _00547_ net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06095_ ci_neuron.uut_simple_neuron.x2\[29\] _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold245 ci_neuron.uut_simple_neuron.titan_id_6\[19\] net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold256 internal_ih.received_byte_count\[6\] net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold267 spi_interface_cvonk.state\[2\] net300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold278 ci_neuron.output_memory\[7\] net311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_113_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_84_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09923_ _00028_ net11 ci_neuron.instruction_i\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold289 ci_neuron.output_memory\[24\] net322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05046_ _00715_ _00731_ net241 _00732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09854_ _00433_ clknet_leaf_122_sys_clock_i ci_neuron.output_memory\[22\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08805_ _04224_ _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06997_ _02612_ _02614_ _02630_ _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09785_ _00364_ clknet_leaf_137_sys_clock_i internal_ih.byte4\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05948_ _01605_ _01606_ _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08736_ _04190_ _04194_ _04195_ _00291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05879_ _01464_ _01483_ _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08667_ spi_interface_cvonk.SCLK_r\[2\] _04125_ _04128_ _04135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07618_ _03159_ _03180_ _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08598_ _03861_ _04072_ _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_119_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07549_ _03162_ _03174_ _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09219_ _04034_ _03809_ _04509_ _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_75_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08435__I1 _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08849__I _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_5_0_sys_clock_i clknet_0_sys_clock_i clknet_4_5_0_sys_clock_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_86_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05885__A1 _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07874__A2 ci_neuron.uut_simple_neuron.titan_id_5\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08823__A1 _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09466__I3 _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05637__A1 _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07149__B _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06920_ ci_neuron.uut_simple_neuron.x3\[20\] _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06851_ _02438_ _02485_ _02486_ _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_128_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06782_ _02364_ _02367_ _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05802_ _01428_ _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09570_ ci_neuron.output_val_internal\[29\] _04771_ _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05733_ _01319_ _01350_ _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08521_ _02091_ _04011_ _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_141_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08452_ _03951_ _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_34_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07403_ _03029_ _03030_ _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05664_ _01328_ _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05595_ _01192_ _01224_ _01228_ _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08383_ net453 _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07334_ _01895_ _02313_ _02905_ _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_116_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout5_I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07265_ _02888_ _02894_ _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_115_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06216_ _01866_ _00165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09004_ _04352_ _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07196_ _02825_ _02746_ _02826_ _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_103_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06147_ _01798_ _01801_ _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_57_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06078_ _01691_ _01724_ _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09906_ _00002_ net10 ci_neuron.address_i\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05029_ _00710_ _00714_ _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_70_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07553__A1 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09837_ _00416_ clknet_leaf_90_sys_clock_i ci_neuron.output_memory\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09768_ _00347_ clknet_leaf_138_sys_clock_i internal_ih.byte2\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08719_ _04177_ _04179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_96_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09699_ net62 clknet_leaf_132_sys_clock_i spi_interface_cvonk.SS_r\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07856__A2 ci_neuron.uut_simple_neuron.titan_id_5\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06652__I _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05380_ ci_neuron.uut_simple_neuron.x2\[14\] _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07050_ _02682_ _02680_ _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06283__A1 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06001_ _01614_ _01615_ _01658_ _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_88_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07607__B ci_neuron.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07952_ net416 _00140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06903_ _02531_ _02537_ _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07883_ net564 net304 _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06834_ _02425_ _02426_ _02429_ _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08583__I0 _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ net332 ci_neuron.output_memory\[14\] _04805_ _04808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09553_ _03935_ _04761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06765_ net40 _02349_ _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_108_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08504_ _03951_ _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06696_ _02283_ _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05716_ _01379_ _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09484_ _04701_ _04702_ _04703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_47_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05647_ _01306_ _01307_ _01312_ _01313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_109_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08435_ ci_neuron.normalised_stream_write_address\[1\] _03935_ _03927_ _03936_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_136_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08366_ ci_neuron.uut_simple_neuron.x0\[24\] _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05578_ _01240_ _01245_ _01246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07317_ _02547_ _02876_ _02875_ _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_74_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07996__C ci_neuron.uut_simple_neuron.titan_id_5\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08297_ net732 net542 _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__09460__A1 ci_neuron.output_memory\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07248_ _02873_ _02877_ _02878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_12_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_131_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07179_ _02617_ _02737_ _02809_ _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09212__A1 _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10190_ net94 clknet_leaf_78_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06577__A2 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08810__I1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07526__A1 _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_83_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09279__A1 _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05068__A2 _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_14_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_8_sys_clock_i clknet_4_4_0_sys_clock_i clknet_leaf_8_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_125_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_04880_ internal_ih.byte7\[7\] _00616_ _00623_ _00597_ _00624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06550_ _01933_ _02049_ _02192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_88_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06481_ _02080_ _02106_ _02123_ _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05501_ _01137_ _01143_ _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05432_ _01099_ _01102_ _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08220_ net511 net212 _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_145_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05363_ _00743_ _01008_ _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08151_ _03688_ net743 _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07102_ _02623_ _02734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05294_ _00863_ _00967_ _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08082_ net560 _00067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_136_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07033_ _01862_ _02665_ _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_113_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06559__A2 _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08984_ _04339_ _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07935_ net723 _00136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07866_ net541 _00156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09605_ net317 _00557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07797_ net594 net648 _03395_ _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06817_ _02181_ _02453_ _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_06748_ _02335_ _02338_ _02385_ _02386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09536_ _03877_ ci_neuron.input_memory\[1\]\[24\] _01475_ _02865_ _04738_ _04739_
+ _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
Xclkbuf_leaf_71_sys_clock_i clknet_4_12_0_sys_clock_i clknet_leaf_71_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_65_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09467_ _04677_ _04687_ _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06679_ _02316_ _02317_ _02318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08418_ net647 net551 _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_81_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09398_ ci_neuron.output_memory\[4\] _04628_ _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08349_ _03856_ _03859_ _03860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_129_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05470__A2 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10242_ _00139_ clknet_leaf_120_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08795__I0 _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10173_ _00070_ clknet_leaf_61_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09018__I internal_ih.data_pointer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09424__A1 ci_neuron.output_memory\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold608 _03373_ net641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_123_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold619 ci_neuron.uut_simple_neuron.titan_id_4\[1\] net652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09578__I2 ci_neuron.uut_simple_neuron.x2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08786__I0 _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05981_ _01637_ _01639_ _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07720_ net456 ci_neuron.uut_simple_neuron.titan_id_3\[13\] _03332_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04932_ _00656_ _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07651_ net652 net408 _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04863_ internal_ih.byte4\[2\] internal_ih.byte3\[2\] _00608_ _00612_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07582_ _03200_ _03207_ _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06602_ _02170_ _02198_ _02242_ _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05516__A3 _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_113_sys_clock_i clknet_4_9_0_sys_clock_i clknet_leaf_113_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06533_ _01926_ _02044_ _02174_ _02175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_105_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09321_ _04064_ net78 _04572_ _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09502__I2 _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06464_ _02075_ _02077_ _02107_ _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_63_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09252_ _04116_ _03915_ _04490_ _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout21_I net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06395_ _01997_ _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05415_ _01084_ _01085_ _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_90_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09183_ _04487_ _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08203_ _03732_ _00193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09415__A1 ci_neuron.output_memory\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05346_ _01002_ _00983_ _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08134_ _03672_ net615 _03675_ _03676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_60_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05277_ _00951_ _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08065_ net724 ci_neuron.uut_simple_neuron.titan_id_0\[10\] _03619_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07016_ _01831_ _02592_ _02649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_116_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08967_ internal_ih.byte7\[1\] net339 _04327_ _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07918_ net800 ci_neuron.uut_simple_neuron.titan_id_5\[15\] _03496_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08898_ net433 _00356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_20_sys_clock_i clknet_4_6_0_sys_clock_i clknet_leaf_20_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_27_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07849_ _03434_ _03435_ _03438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_84_sys_clock_i_I clknet_4_14_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09519_ _04721_ _04729_ _04731_ _04732_ _00537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__08457__A2 _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_104_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_78_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10225_ _00152_ clknet_leaf_90_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08788__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10156_ _00221_ clknet_leaf_35_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[30\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10087_ _00184_ clknet_leaf_12_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05200_ _00854_ _00874_ _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09248__I1 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06180_ _01832_ _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05131_ ci_neuron.uut_simple_neuron.x2\[6\] _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold427 _03535_ net460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold416 internal_ih.byte5\[2\] net449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_20_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold405 _04320_ net438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05062_ _00746_ _00159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold449 internal_ih.byte3\[6\] net482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold438 ci_neuron.stream_o\[21\] net471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09870_ _00061_ net29 ci_neuron.value_i\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08821_ _04099_ _04237_ _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05964_ _01621_ _01622_ _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08752_ _04194_ net268 _00297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_hold270_I ci_neuron.stream_o\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07703_ _03313_ _03316_ _03318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_04915_ _00639_ _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08683_ _04134_ net126 _04150_ _00283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07634_ _03010_ _03248_ _03258_ _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_05895_ _01520_ _01543_ _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06698__A1 _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04846_ _00596_ _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07565_ _03190_ _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07496_ _03121_ _03122_ _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06516_ net53 _02111_ _02159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06745__I ci_neuron.uut_simple_neuron.x3\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09304_ _04023_ net96 _04561_ _04563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06447_ _02090_ _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09235_ _04074_ _03851_ _04519_ _04521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06378_ _01943_ _01979_ _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09166_ _04479_ _00437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05329_ _00970_ _00940_ _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08117_ _03660_ _03661_ _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09097_ _04417_ ci_neuron.stream_o\[6\] ci_neuron.stream_o\[22\] _04418_ _04438_
+ _04439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_08048_ net603 ci_neuron.uut_simple_neuron.titan_id_0\[7\] ci_neuron.uut_simple_neuron.titan_id_1\[6\]
+ ci_neuron.uut_simple_neuron.titan_id_0\[6\] _03604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_clkbuf_leaf_72_sys_clock_i_I clknet_4_12_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10010_ net76 clknet_leaf_68_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09999_ _00514_ clknet_leaf_103_sys_clock_i internal_ih.expected_byte_count\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05361__A1 _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08602__A2 _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_141_sys_clock_i_I clknet_4_0_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07169__A2 ci_neuron.uut_simple_neuron.x3\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10208_ _00104_ clknet_leaf_119_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10139_ _00204_ clknet_leaf_55_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04927__B2 internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07341__A2 _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05680_ _00740_ _01344_ _01329_ _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__05352__A1 _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07350_ _02916_ _02978_ _02979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06301_ _01935_ _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07281_ _02784_ _02833_ _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05104__A1 _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08841__A2 _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09020_ ci_neuron.output_val_internal\[24\] ci_neuron.output_val_internal\[16\] ci_neuron.output_val_internal\[8\]
+ ci_neuron.output_val_internal\[0\] _04366_ _04367_ _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06232_ _01829_ _01881_ _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_115_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08780__I _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06163_ _01807_ _01815_ _01817_ _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_53_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold202 net699 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05114_ _00793_ _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold213 ci_neuron.uut_simple_neuron.titan_id_6\[9\] net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold235 _04205_ net268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold224 ci_neuron.uut_simple_neuron.titan_id_6\[22\] net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06094_ _01714_ _01715_ _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold257 _04203_ net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold246 internal_ih.current_instruction\[0\] net279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold268 _04541_ net301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_113_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09922_ _00027_ net11 ci_neuron.instruction_i\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xhold279 _04799_ net312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05045_ _00728_ _00730_ _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09853_ _00432_ clknet_leaf_120_sys_clock_i ci_neuron.output_memory\[21\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08804_ net275 _04236_ _04238_ _00316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09784_ _00363_ clknet_leaf_145_sys_clock_i internal_ih.byte4\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06996_ _02619_ _02627_ _02629_ _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_08735_ net256 _04189_ _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05947_ _01567_ _01588_ _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05878_ _01464_ _01483_ _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08666_ _04133_ _04134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_37_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07617_ _03240_ _03241_ _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08597_ _03862_ _04072_ _04076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07548_ _03172_ _03173_ _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_60_sys_clock_i_I clknet_4_15_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07479_ _03105_ _03106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_118_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09218_ _04511_ _00457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09149_ net218 _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold780 _01961_ net824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__04909__A1 internal_ih.byte5\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_19_sys_clock_i_I clknet_4_6_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08823__A2 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08533__C _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08587__A1 ci_neuron.value_i\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06850_ _02440_ _02456_ _02486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05801_ _01428_ _01431_ _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08976__S _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06781_ _02359_ _02416_ _02417_ _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_128_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05732_ _00932_ _01395_ _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08775__I _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08520_ _03939_ _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10022__D net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05663_ _01327_ _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08511__A1 _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08451_ _03950_ _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_34_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07402_ _01969_ _02957_ _03030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05594_ _01083_ _01210_ _01176_ _01260_ _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_58_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08382_ net331 _00186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07333_ _02961_ _02922_ _02962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_128_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07264_ _02891_ _02893_ _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06215_ _01851_ _01865_ _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_60_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09003_ _04173_ _04174_ _04181_ _04192_ _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_07195_ _02276_ _02745_ _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06146_ _01699_ _01799_ _01800_ _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_57_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06077_ _01733_ _00220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_70_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09905_ _00024_ net12 ci_neuron.address_i\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05028_ ci_neuron.instruction_i\[0\] ci_neuron.instruction_i\[1\] _00713_ _00714_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_70_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09836_ _00415_ clknet_leaf_89_sys_clock_i ci_neuron.output_memory\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06979_ _02550_ _02559_ _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09767_ _00346_ clknet_leaf_127_sys_clock_i internal_ih.byte2\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09698_ net2 clknet_leaf_133_sys_clock_i spi_interface_cvonk.SS_r\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08718_ net313 _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05316__A1 _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08502__A1 _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08649_ _04119_ net531 _04111_ _04120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_68_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09302__I0 _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_7_sys_clock_i clknet_4_4_0_sys_clock_i clknet_leaf_7_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07480__A1 _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06000_ _01580_ _01613_ _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_70_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_110_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07951_ _03522_ net415 _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06902_ _02536_ _02534_ _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_120_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07882_ net306 _00158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_52_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06833_ _02469_ _00237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08583__I1 _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09621_ net372 _00564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06764_ net40 _02349_ _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09552_ _03930_ _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_108_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05715_ ci_neuron.uut_simple_neuron.x2\[21\] ci_neuron.uut_simple_neuron.x2\[22\]
+ _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08503_ _03986_ _03994_ _03995_ _00258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09288__A2 _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06695_ _02283_ _02333_ _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_78_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70_sys_clock_i clknet_4_12_0_sys_clock_i clknet_leaf_70_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09483_ _03822_ ci_neuron.input_memory\[1\]\[16\] _01150_ _02384_ _04691_ _04692_
+ _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_47_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05646_ _01309_ _01277_ _01311_ _01312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_93_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08434_ ci_neuron.address_i\[1\] _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_135_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05577_ _01243_ _01244_ _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08365_ _03873_ _00184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07316_ _02926_ _02944_ _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08296_ _03813_ _00175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06274__A2 _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07247_ _02547_ _02876_ _02877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07178_ _02808_ _02736_ _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09212__A2 _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06129_ _01743_ _01775_ _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06329__A3 _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09819_ _00398_ clknet_leaf_134_sys_clock_i internal_ih.current_instruction\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_89_sys_clock_i clknet_4_11_0_sys_clock_i clknet_leaf_89_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_127_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07462__A1 _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07214__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09214__I _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_112_sys_clock_i clknet_4_10_0_sys_clock_i clknet_leaf_112_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06480_ _02084_ _02105_ _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05500_ _01130_ _01167_ _01168_ _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_74_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05431_ _01100_ _01101_ _00963_ _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_83_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08150_ net742 net811 _03689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07101_ _02620_ _02681_ _02732_ _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05362_ _00888_ _00985_ _01033_ _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_83_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05293_ _00891_ _00914_ _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08081_ _03631_ _03632_ _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_136_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07032_ _02175_ _02193_ _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold398_I internal_ih.byte4\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08983_ _04339_ _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07934_ _03508_ net722 _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07865_ net540 _03451_ _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_hold732_I _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09604_ ci_neuron.stream_o\[6\] net316 _04795_ _04798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07796_ _03387_ _03388_ _03394_ _03391_ _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06816_ _02144_ _02285_ _02453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_06747_ _02333_ _02384_ _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09535_ _04700_ _04746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06678_ _01891_ _01938_ _02317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09466_ _03809_ ci_neuron.input_memory\[1\]\[14\] _01052_ _02335_ _04667_ _04669_
+ _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_65_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05629_ _01288_ _01294_ _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08417_ _03917_ _03918_ _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09397_ _04599_ _04628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08348_ _03844_ _03846_ _03857_ _03858_ _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_19_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08279_ _03795_ _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05099__I _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10241_ _00137_ clknet_leaf_120_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08795__I1 _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10172_ _00069_ clknet_leaf_60_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_38_sys_clock_i clknet_4_5_0_sys_clock_i clknet_leaf_38_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_85_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold609 ci_neuron.uut_simple_neuron.titan_id_1\[23\] net642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_52_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09188__A1 _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05980_ _01597_ _01598_ _01638_ _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04931_ internal_ih.byte6\[2\] _00652_ _00653_ internal_ih.byte2\[2\] _00656_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07650_ _03274_ _00249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04862_ _00611_ _00026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07581_ _01833_ _03206_ _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06601_ _02172_ _02197_ _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06532_ _02173_ _02148_ _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09320_ _04566_ _04572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_48_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09502__I3 _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09251_ _04529_ _00472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_138_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06463_ _02080_ _02106_ _02107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_91_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08202_ _03726_ _03730_ _03731_ _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06394_ _01867_ _02038_ _02039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05414_ _01047_ _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09182_ _04488_ _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05345_ _01017_ _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08133_ net614 ci_neuron.uut_simple_neuron.titan_id_0\[21\] _03675_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_60_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08064_ _03614_ _03616_ _03617_ _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_4_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07015_ _02639_ _02637_ _02647_ _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_114_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05276_ _00931_ _00933_ _00950_ _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_70_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08966_ net344 _00386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07917_ ci_neuron.uut_simple_neuron.titan_id_2\[15\] ci_neuron.uut_simple_neuron.titan_id_5\[15\]
+ _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08897_ internal_ih.byte3\[2\] net432 _04291_ _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07848_ ci_neuron.uut_simple_neuron.titan_id_2\[4\] net590 _03437_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07779_ net611 _03380_ _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09518_ net188 _04727_ _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09873__CLK net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09449_ _04649_ _04665_ _04671_ _04672_ _00527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_132_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10224_ _00149_ clknet_leaf_93_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10155_ _00220_ clknet_leaf_35_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08868__I _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10086_ _00183_ clknet_leaf_12_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08940__I1 internal_ih.byte4\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07408__A1 _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05130_ _00808_ _00809_ _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07959__A2 net458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_133_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08081__A1 _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold406 internal_ih.byte5\[3\] net439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold417 _04323_ net450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__04890__B2 internal_ih.byte0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05061_ _00737_ _00745_ _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold439 _04818_ net472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold428 _03537_ net461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09746__CLK clknet_4_4_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08820_ _04247_ _00323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05963_ ci_neuron.uut_simple_neuron.x2\[1\] ci_neuron.uut_simple_neuron.x2\[27\]
+ _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08751_ net267 _04204_ _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05894_ _01520_ _01543_ _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07702_ net413 _00126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04914_ _00645_ _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08682_ _04146_ _04149_ _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07633_ _03251_ _03254_ _03257_ _03258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_49_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04845_ internal_ih.current_instruction\[3\] _00592_ _00593_ _00595_ _00596_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_71_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07564_ _03187_ _03189_ _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_119_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09097__B1 ci_neuron.stream_o\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09402__I _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07495_ _03031_ _03037_ _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06515_ _02154_ _02157_ _02158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_76_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09303_ _04562_ _00491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_62_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06446_ ci_neuron.uut_simple_neuron.x3\[10\] _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09234_ _04520_ _00464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09165_ net99 _04479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06377_ _02016_ _02022_ _02023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08116_ _03657_ net584 _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05328_ _00892_ _01000_ _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09096_ _04405_ _04437_ _04438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05259_ _00905_ _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08047_ _03594_ _03599_ _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09411__I2 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09572__A1 ci_neuron.output_memory\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__A1 _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09998_ net159 clknet_leaf_102_sys_clock_i internal_ih.expected_byte_count\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08949_ net339 net403 _04317_ _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06310__A1 _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05287__I _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10207_ _00103_ clknet_leaf_48_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10138_ _00203_ clknet_leaf_56_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10069_ _00196_ clknet_leaf_82_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08547__B _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05750__I _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07280_ _02847_ _02850_ _02909_ _02910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_06300_ _01946_ _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06231_ net37 _01877_ _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_116_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06162_ _01779_ _01781_ _01816_ _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06093_ _01747_ _01748_ _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05113_ _00756_ _00766_ _00793_ _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
Xhold203 _04443_ net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold214 ci_neuron.uut_simple_neuron.titan_id_6\[3\] net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold225 ci_neuron.output_val_internal\[30\] net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_111_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold258 ci_neuron.uut_simple_neuron.x0\[22\] net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold247 _00394_ net280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold269 _00479_ net302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold236 internal_ih.byte2\[3\] net269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09921_ _00026_ net21 ci_neuron.instruction_i\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05044_ _00708_ _00729_ _00713_ _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_41_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__A1 _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_123_Left_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09852_ _00431_ clknet_leaf_120_sys_clock_i ci_neuron.output_memory\[20\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08803_ _04059_ _04237_ _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09783_ _00362_ clknet_leaf_144_sys_clock_i internal_ih.byte4\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06995_ _02329_ _02628_ _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08734_ _04193_ _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05946_ _01572_ _01587_ _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05877_ _01523_ _01537_ _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08665_ _04124_ _04133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07616_ _02550_ _03178_ _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08596_ _04075_ _00271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_132_Left_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07547_ _02733_ _02736_ _03012_ _03173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_49_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07478_ _03078_ _03104_ _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06429_ _02013_ _02031_ net54 _02062_ _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_106_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09217_ _04027_ _03797_ _04509_ _04511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09911__CLK net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09148_ _04470_ _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09079_ ci_neuron.output_val_internal\[28\] ci_neuron.output_val_internal\[20\] ci_neuron.output_val_internal\[12\]
+ ci_neuron.output_val_internal\[4\] _04390_ _04391_ _04423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_130_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_141_Left_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_130_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_6_sys_clock_i clknet_4_4_0_sys_clock_i clknet_leaf_6_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold770 internal_ih.byte1\[4\] net814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold781 ci_neuron.uut_simple_neuron.titan_id_2\[23\] net825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07020__A2 _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05334__A2 _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08587__A2 _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08831__I0 _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05270__A1 _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05800_ _01461_ _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06780_ _02361_ _02400_ _02417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_128_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05731_ _01359_ _01394_ _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07314__A3 _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05662_ _01326_ _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08450_ _03934_ _03950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_34_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07401_ _02374_ _02395_ _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08381_ _03886_ net330 _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07332_ _02950_ _02960_ _02961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05593_ _00887_ _01210_ _01211_ _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_86_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07078__A2 _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07263_ _01935_ _02892_ _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07194_ _02225_ _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06214_ _01857_ _01864_ _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09002_ _04350_ _04254_ _04178_ _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06145_ _01746_ _01770_ _01699_ _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06589__A1 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06076_ _01729_ _01732_ _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09904_ _00023_ net12 ci_neuron.address_i\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05027_ ci_neuron.instruction_i\[2\] _00711_ _00712_ _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA_hold762_I internal_ih.byte1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09835_ _00414_ clknet_leaf_90_sys_clock_i ci_neuron.output_memory\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06978_ _02178_ _02611_ _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09766_ _00345_ clknet_leaf_127_sys_clock_i internal_ih.byte1\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05929_ _01568_ _01588_ _01589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08717_ _04173_ _04176_ net313 _04177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09697_ net770 clknet_leaf_132_sys_clock_i spi_interface_cvonk.SCLK_r\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_88_sys_clock_i clknet_4_11_0_sys_clock_i clknet_leaf_88_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08648_ ci_neuron.value_i\[30\] _04118_ _04026_ _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_68_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08579_ _03840_ _04044_ _03852_ _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_49_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05004__A1 internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06752__A1 _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_111_sys_clock_i clknet_4_10_0_sys_clock_i clknet_leaf_111_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06396__I _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_123_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09500__I _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07480__A2 _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05491__A1 _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07950_ ci_neuron.uut_simple_neuron.titan_id_2\[21\] net414 _03523_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06901_ _02535_ _01832_ _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07881_ net305 _03465_ _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_52_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06832_ _02466_ _02468_ _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09620_ net371 ci_neuron.output_memory\[13\] _04805_ _04807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06763_ _02359_ _02361_ _02400_ _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09551_ ci_neuron.output_memory\[27\] _04744_ _04759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_108_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05714_ _01146_ _01376_ _01377_ _01378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08502_ _01998_ _03980_ _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06694_ ci_neuron.uut_simple_neuron.x3\[15\] _02333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09482_ _04700_ _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_47_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05645_ _01279_ _01310_ _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08433_ _03929_ _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05576_ _01123_ _01162_ _01200_ _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_117_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08364_ _03869_ _03872_ _03873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07315_ _02942_ _02943_ _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_73_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08295_ _03809_ _03810_ _03812_ _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_6_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07246_ _02874_ _02875_ _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07177_ _02726_ _02806_ _02807_ _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_5_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06128_ _01771_ _01774_ _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06059_ _01714_ _01715_ _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xclkbuf_leaf_37_sys_clock_i clknet_4_5_0_sys_clock_i clknet_leaf_37_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09818_ _00397_ clknet_leaf_132_sys_clock_i internal_ih.current_instruction\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_97_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09749_ _00328_ clknet_leaf_33_sys_clock_i ci_neuron.uut_simple_neuron.x2\[30\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08629__C _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_83_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09320__I _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05473__A1 _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09054__I3 ci_neuron.output_val_internal\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05225__A1 _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05430_ _00969_ _01005_ ci_neuron.uut_simple_neuron.x2\[14\] _01101_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_74_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05361_ _01012_ _01020_ _01033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07100_ _02623_ _02731_ _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_56_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05292_ _00941_ _00943_ _00965_ _00916_ _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_08080_ net518 net559 _03632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07031_ _02662_ _02611_ _02663_ _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09045__I3 ci_neuron.output_val_internal\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05216__A1 ci_neuron.uut_simple_neuron.x2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_143_Right_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08982_ _04183_ _04185_ _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07933_ net721 ci_neuron.uut_simple_neuron.titan_id_5\[18\] _03509_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_138_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07864_ ci_neuron.uut_simple_neuron.titan_id_2\[7\] ci_neuron.uut_simple_neuron.titan_id_5\[7\]
+ _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_hold460_I internal_ih.byte2\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06815_ _02444_ _02451_ _02452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_3_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09603_ net308 _00556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07795_ net594 ci_neuron.uut_simple_neuron.titan_id_3\[26\] _03394_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06746_ _02383_ _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_79_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold725_I _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09534_ ci_neuron.output_memory\[24\] _04744_ _04745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06677_ _01891_ _01938_ _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_94_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09465_ ci_neuron.output_memory\[14\] _04675_ _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_109_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05628_ _01292_ _01293_ _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08416_ _03910_ _03913_ _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_22_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09396_ _04597_ _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05559_ _01226_ _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08347_ _03836_ _03850_ net390 _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08278_ _03795_ _03797_ _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08641__A1 _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07229_ _02801_ _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10240_ _00136_ clknet_leaf_115_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10171_ _00068_ clknet_leaf_60_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_68_sys_clock_i_I clknet_4_12_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09188__A2 _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04930_ _00655_ _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_0_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04861_ internal_ih.byte7\[1\] _00606_ _00609_ _00610_ _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06600_ _02213_ _02215_ _02240_ _02241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07580_ _03203_ _03205_ _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06531_ _01925_ _02173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_105_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07123__A1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09250_ _04110_ _03904_ _04525_ _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_138_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06462_ _02084_ _02105_ _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08201_ _03724_ _03727_ _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06393_ _01853_ _01925_ _02037_ _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05413_ _01044_ _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09181_ _04487_ _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05344_ _00976_ _01015_ _01016_ _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_60_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08132_ net616 _00076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_137_sys_clock_i_I clknet_4_0_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05275_ _00934_ _00949_ _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08063_ net561 ci_neuron.uut_simple_neuron.titan_id_0\[9\] net654 ci_neuron.uut_simple_neuron.titan_id_0\[8\]
+ _03617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07014_ _02634_ _02636_ _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_101_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08965_ net343 internal_ih.byte6\[0\] _04327_ _04330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07916_ net748 _00133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08896_ _04290_ _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09351__A2 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07847_ net737 _00153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07778_ _03376_ _03377_ _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10221__D _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06729_ _02366_ _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09517_ _04724_ _04730_ _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09448_ net103 _04655_ _04672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09379_ ci_neuron.output_memory\[1\] _04600_ _04613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_7_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_18_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10223_ _00138_ clknet_leaf_93_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10154_ _00219_ clknet_leaf_36_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10085_ _00182_ clknet_leaf_19_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_56_sys_clock_i_I clknet_4_15_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold418 internal_ih.spi_rx_byte_i\[4\] net451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold407 _04314_ net440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05060_ _00744_ _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold429 internal_ih.byte3\[5\] net462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_36_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06919__A1 _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05962_ _01618_ _01620_ _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08750_ internal_ih.received_byte_count\[6\] _04202_ _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07344__A1 _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05893_ _01553_ _00216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07701_ net412 _03316_ _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_04913_ internal_ih.byte5\[3\] _00640_ _00641_ internal_ih.byte1\[3\] _00645_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08681_ _04148_ _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_125_sys_clock_i_I clknet_4_3_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07632_ _03255_ _03256_ _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_49_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04844_ _00594_ internal_ih.current_instruction\[2\] _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_45_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07563_ _02132_ _03188_ _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09302_ _04017_ net84 _04561_ _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07494_ _03034_ _03036_ _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06514_ _02075_ _02155_ _02156_ _02157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06445_ _02001_ _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09233_ _04069_ _03849_ _04519_ _04520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09164_ _04478_ _00436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06376_ _02017_ _02020_ _02021_ _02022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08115_ net583 net670 _03660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05327_ _00886_ _00914_ _00984_ _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09095_ _04419_ ci_neuron.stream_o\[14\] _04437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05258_ _00932_ _00921_ _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08046_ _03588_ _03591_ _03601_ _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_4_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05189_ net675 _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08969__I _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_5_sys_clock_i clknet_4_1_0_sys_clock_i clknet_leaf_5_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_73_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09411__I3 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07583__A1 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09997_ _00512_ clknet_leaf_102_sys_clock_i internal_ih.expected_byte_count\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08948_ net438 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08879_ _04281_ _00348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05568__I _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_44_sys_clock_i_I clknet_4_7_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05821__A1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10206_ _00102_ clknet_leaf_48_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09563__A2 _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10137_ _00202_ clknet_leaf_55_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10068_ _00195_ clknet_leaf_80_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07326__A1 _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06230_ _01838_ _01879_ _01880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06161_ _01737_ _01778_ _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06092_ _01663_ _01717_ _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05112_ ci_neuron.uut_simple_neuron.x2\[5\] _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold204 ci_neuron.uut_simple_neuron.titan_id_6\[29\] net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold226 _00546_ net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_leaf_113_sys_clock_i_I clknet_4_9_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold215 ci_neuron.uut_simple_neuron.titan_id_6\[7\] net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_123_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05812__A1 _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold259 _03861_ net292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold248 internal_ih.current_instruction\[5\] net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold237 _04293_ net270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09920_ _00025_ net20 ci_neuron.instruction_i\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05043_ _00709_ _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_113_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09851_ _00430_ clknet_leaf_115_sys_clock_i ci_neuron.output_memory\[19\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06994_ net49 _02447_ _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08802_ _04207_ _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09782_ _00361_ clknet_leaf_145_sys_clock_i internal_ih.byte3\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05945_ _01602_ _01603_ _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08733_ _04191_ _04192_ _04187_ _04188_ _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
Xclkbuf_leaf_87_sys_clock_i clknet_4_11_0_sys_clock_i clknet_leaf_87_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05876_ _01527_ _01536_ _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08664_ _04130_ net254 _00282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_37_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07615_ _02559_ _03177_ _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08595_ _04074_ _02804_ _04053_ _04075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07546_ _03165_ _03171_ _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07477_ _03100_ _03103_ _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09216_ _04510_ _00456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06428_ _02029_ _02071_ _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06359_ _01926_ _02004_ _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09147_ net146 _04470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06056__A1 _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09078_ _04417_ ci_neuron.stream_o\[4\] ci_neuron.stream_o\[20\] _04418_ _04421_
+ _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_32_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08029_ _03584_ _03586_ _03587_ _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xhold760 ci_neuron.uut_simple_neuron.titan_id_0\[25\] net811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_12_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold771 internal_ih.byte1\[2\] net815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold782 ci_neuron.uut_simple_neuron.titan_id_5\[29\] net826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07556__A1 _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_13_0_sys_clock_i clknet_0_sys_clock_i clknet_4_13_0_sys_clock_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_110_sys_clock_i clknet_4_8_0_sys_clock_i clknet_leaf_110_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_32_sys_clock_i_I clknet_4_4_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07547__A1 _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08595__I0 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_129_sys_clock_i clknet_4_2_0_sys_clock_i clknet_leaf_129_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_128_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05730_ _01361_ _01366_ _01393_ _01394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_89_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05661_ _01266_ _01290_ _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_101_sys_clock_i_I clknet_4_8_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07400_ _03027_ _03001_ _03028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08380_ net329 net396 _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_34_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07331_ _02953_ _02959_ _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_128_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05592_ _01221_ _01230_ _01258_ _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07262_ _02323_ _02344_ _02892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_128_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07193_ _02822_ _02823_ _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06213_ _01863_ _01864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09001_ net26 _04350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06144_ _01746_ _01770_ _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_112_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06075_ _01730_ _01731_ _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09903_ _00022_ net12 ci_neuron.address_i\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05026_ ci_neuron.instruction_i\[4\] ci_neuron.instruction_i\[7\] ci_neuron.instruction_i\[6\]
+ _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xclkbuf_leaf_36_sys_clock_i clknet_4_5_0_sys_clock_i clknet_leaf_36_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_70_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09834_ _00413_ clknet_4_11_0_sys_clock_i ci_neuron.output_memory\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06210__A1 _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06977_ _02610_ _02146_ _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_09765_ _00344_ clknet_leaf_127_sys_clock_i internal_ih.byte1\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xrebuffer30 _02142_ net500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05928_ _01572_ _01587_ _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09696_ net63 clknet_leaf_132_sys_clock_i spi_interface_cvonk.SCLK_r\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08716_ _04174_ _04175_ _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_139_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05859_ _01467_ _01486_ _01519_ _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_96_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08647_ _03916_ _03910_ _04107_ _04118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_68_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08578_ _04060_ _00268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07529_ _03154_ _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_119_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_81_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold590 _03585_ net623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08577__I0 _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_20_sys_clock_i_I clknet_4_6_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09254__S _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05555__A3 _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06504__A2 _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_123_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06900_ _02102_ _02079_ _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07880_ ci_neuron.uut_simple_neuron.titan_id_2\[9\] ci_neuron.uut_simple_neuron.titan_id_5\[9\]
+ _03465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_52_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06831_ _02467_ _02406_ _02410_ _02414_ _02468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_06762_ _02369_ _02399_ _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09550_ _04743_ _04755_ _04757_ _04758_ _00542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_37_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05713_ _01375_ _01336_ _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08501_ ci_neuron.value_i\[8\] _03944_ _03993_ _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_37_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09481_ _00728_ _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06693_ _02182_ net50 _02331_ _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_108_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08432_ _03928_ _03932_ _03933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08496__A2 _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05644_ _01247_ _01308_ _01277_ _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_93_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05575_ _01242_ _01241_ _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08363_ _03866_ _03870_ _03871_ _03865_ _03872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_144_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07314_ _02554_ _02557_ _02733_ _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08294_ _03803_ _03806_ _03811_ _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07245_ _02548_ _02680_ _02875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07176_ _02804_ _02805_ _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06127_ _01782_ _00221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06431__A1 _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06058_ ci_neuron.uut_simple_neuron.x2\[29\] _01670_ _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05009_ _00700_ _00052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09817_ _00396_ clknet_leaf_133_sys_clock_i internal_ih.current_instruction\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09748_ _00327_ clknet_leaf_33_sys_clock_i ci_neuron.uut_simple_neuron.x2\[29\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06498__A1 _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09679_ _00266_ clknet_leaf_48_sys_clock_i ci_neuron.uut_simple_neuron.x3\[16\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05170__A1 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09436__A1 ci_neuron.output_memory\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04984__A1 internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_3_sys_clock_i_I clknet_4_1_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05360_ _01001_ _01030_ _01031_ _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05291_ _00739_ _00964_ _00965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07030_ _02146_ _02610_ _02663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08981_ net374 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07932_ ci_neuron.uut_simple_neuron.titan_id_2\[17\] ci_neuron.uut_simple_neuron.titan_id_5\[17\]
+ _03497_ _03505_ _03507_ _03508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_07863_ ci_neuron.uut_simple_neuron.titan_id_2\[6\] net539 _03449_ _03450_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06814_ _02330_ _02450_ _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_74_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08961__I0 internal_ih.byte6\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09602_ ci_neuron.stream_o\[5\] net307 _04795_ _04797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07794_ _03393_ _00113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09533_ _04674_ _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06745_ ci_neuron.uut_simple_neuron.x3\[16\] _02383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06676_ _02312_ _02314_ _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09464_ _04673_ _04682_ _04684_ _04685_ _00529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05627_ _01263_ _01267_ _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_80_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08415_ _03915_ _03916_ _03917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09395_ _04598_ _04621_ _04625_ _04626_ _00519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_08346_ net390 net429 _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_22_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05558_ ci_neuron.uut_simple_neuron.x2\[18\] _01226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05489_ _01081_ _01113_ _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08277_ _03796_ _03797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10219__D _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07228_ _02799_ _02858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07159_ _02720_ _02748_ _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_104_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06404__A1 _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ _00067_ clknet_leaf_59_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08952__I0 internal_ih.byte6\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09106__B1 ci_neuron.stream_o\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06955__I _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09331__I _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_127_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08632__A2 _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09506__I _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04860_ _00596_ _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06530_ _02134_ _02150_ _02171_ _02172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_105_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06461_ _02099_ _02104_ _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_138_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05412_ _00887_ _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08200_ _03729_ _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06392_ _01852_ _02007_ _02037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09180_ _04486_ _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05343_ _01013_ _01014_ _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_83_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08131_ _03672_ net615 _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_60_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08623__A2 _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06634__A1 _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05274_ _00935_ _00948_ _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08062_ _03606_ _03615_ _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07013_ _02646_ _00240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_4_sys_clock_i clknet_4_1_0_sys_clock_i clknet_leaf_4_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_141_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08964_ net346 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07915_ net747 ci_neuron.uut_simple_neuron.titan_id_5\[15\] _03493_ _03494_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09416__I _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08895_ _04256_ _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09351__A3 _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07846_ net736 _03435_ _03436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07777_ ci_neuron.uut_simple_neuron.titan_id_4\[23\] net610 _03379_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04989_ _00689_ _00042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06728_ _01947_ _01988_ _02365_ _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09516_ _03851_ ci_neuron.input_memory\[1\]\[21\] _01368_ _02804_ _04716_ _04717_
+ _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_39_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09447_ _04652_ _04670_ _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06659_ _02259_ _02298_ _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_94_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09378_ _04598_ _04601_ _04609_ _04612_ _00516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_90_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08329_ _03839_ _03842_ _03843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_61_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10222_ _00127_ clknet_leaf_94_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_6\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10153_ _00218_ clknet_leaf_40_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04939__A1 internal_ih.byte6\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05600__A2 _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10084_ _00181_ clknet_leaf_19_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_89_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07105__A2 _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold408 internal_ih.byte0\[3\] net441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_40_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold419 _04262_ net452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07700_ ci_neuron.uut_simple_neuron.titan_id_4\[10\] ci_neuron.uut_simple_neuron.titan_id_3\[10\]
+ _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05961_ _01619_ _01531_ _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05892_ _01550_ _01552_ _01553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_86_sys_clock_i clknet_4_14_0_sys_clock_i clknet_leaf_86_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_04912_ _00644_ _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08680_ _04135_ _04141_ _04147_ _04148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07631_ _02132_ _03188_ _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04843_ net733 _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_144_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07562_ _02542_ _02562_ _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_49_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06513_ _02077_ _02107_ _02156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09301_ _04545_ _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09341__I0 _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07493_ _02898_ _03050_ _03119_ _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_119_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06444_ _01955_ _02052_ _02087_ _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_61_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09232_ _04499_ _04519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_8_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06375_ _02018_ _02019_ _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_32_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09163_ net101 _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05326_ _00997_ _00998_ _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08114_ net585 _00073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09094_ _04415_ net224 _04436_ _00408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_142_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05257_ _00905_ _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_hold785_I _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08045_ ci_neuron.uut_simple_neuron.titan_id_1\[5\] ci_neuron.uut_simple_neuron.titan_id_0\[5\]
+ _03601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_101_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05188_ ci_neuron.uut_simple_neuron.x2\[6\] _00861_ _00866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_73_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09996_ _00511_ clknet_leaf_11_sys_clock_i ci_neuron.input_memory\[1\]\[31\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08947_ net437 internal_ih.byte5\[0\] _04317_ _04320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08878_ net432 net481 _04280_ _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07829_ net567 ci_neuron.uut_simple_neuron.titan_id_5\[1\] _03422_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_98_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09332__I0 _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05821__A2 _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07023__A1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10205_ _00101_ clknet_leaf_61_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10136_ _00201_ clknet_leaf_55_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_128_sys_clock_i clknet_4_3_0_sys_clock_i clknet_leaf_128_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10067_ _00194_ clknet_leaf_79_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09323__I0 _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06160_ _01767_ _01809_ _01814_ _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_81_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07262__A1 _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06091_ _01707_ _01708_ _01716_ _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05111_ _00791_ _00767_ _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold205 internal_ih.spi_tx_byte_o\[3\] net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold216 spi_interface_cvonk.state\[1\] net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold227 ci_neuron.uut_simple_neuron.x2\[26\] net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold249 internal_ih.current_instruction\[6\] net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold238 internal_ih.received_byte_count\[3\] net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_22_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05042_ _00727_ _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_40_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_35_sys_clock_i clknet_4_5_0_sys_clock_i clknet_leaf_35_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08762__A1 _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_2_0_sys_clock_i clknet_0_sys_clock_i clknet_4_2_0_sys_clock_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09850_ _00429_ clknet_leaf_114_sys_clock_i ci_neuron.output_memory\[18\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05576__A1 _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06993_ _02495_ _02626_ _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08801_ _04208_ _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09781_ _00360_ clknet_leaf_145_sys_clock_i internal_ih.byte3\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05944_ _01255_ _01566_ _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08732_ _04185_ _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_0_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09562__I0 _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08663_ net253 _04131_ _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05875_ _01535_ _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07614_ ci_neuron.uut_simple_neuron.x3\[30\] _02611_ _03238_ _03239_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09314__I0 _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08594_ _04019_ _04071_ _04072_ _04073_ _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_49_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_138_Right_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07545_ _02939_ _03170_ _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08817__A2 _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07476_ _02497_ _03102_ _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_48_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06427_ _02033_ _02063_ _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09215_ _04023_ _03795_ _04509_ _04510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06358_ _02003_ _02000_ _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09146_ _04469_ _00427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07253__A1 _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06289_ _01824_ _01936_ _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05309_ _00982_ _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06056__A2 _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09077_ _04405_ _04420_ _04421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08028_ ci_neuron.uut_simple_neuron.titan_id_1\[4\] ci_neuron.uut_simple_neuron.titan_id_0\[4\]
+ _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold750 _03397_ net783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold761 ci_neuron.uut_simple_neuron.titan_id_5\[28\] net812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold772 ci_neuron.uut_simple_neuron.titan_id_2\[29\] net816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__05567__A1 _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09979_ _00494_ clknet_leaf_48_sys_clock_i ci_neuron.input_memory\[1\]\[14\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08595__I1 _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10119_ _00243_ clknet_leaf_37_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_128_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05660_ _00859_ _01178_ _01324_ _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_05591_ _01222_ _01229_ _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_34_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07330_ _02956_ _02958_ _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_133_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07483__A1 _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07261_ _02889_ _02818_ _02890_ _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_73_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09000_ _04349_ _00401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07192_ _01883_ _02755_ _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06212_ _01862_ _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06143_ _01749_ _01768_ _01797_ _01798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06074_ _01647_ _01685_ _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_111_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09902_ _00021_ net12 ci_neuron.address_i\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05025_ ci_neuron.instruction_i\[3\] ci_neuron.instruction_i\[5\] _00711_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_hold483_I internal_ih.byte5\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09833_ _00412_ clknet_leaf_93_sys_clock_i ci_neuron.output_memory\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06976_ _02279_ _02561_ _02609_ _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09764_ _00343_ clknet_leaf_134_sys_clock_i internal_ih.byte1\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xrebuffer20 _02108_ net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05927_ _01527_ _01586_ _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09695_ net1 clknet_leaf_133_sys_clock_i spi_interface_cvonk.SCLK_r\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08715_ internal_ih.spi_rx_byte_i\[3\] _04171_ _04175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05858_ _01470_ _01485_ _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08646_ _04117_ _00279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_138_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05789_ _01450_ _01443_ _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05721__A1 _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08577_ _04059_ _02616_ _04053_ _04060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07528_ _03118_ _03132_ _03153_ _03154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07459_ _02934_ _03008_ _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09129_ net264 _04461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold580 net816 net613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold591 ci_neuron.uut_simple_neuron.titan_id_5\[24\] net624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08577__I1 _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06179__B _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_72_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_123_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_81_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07029__I _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06830_ _02256_ _02299_ _02354_ _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06761_ _02372_ _02398_ _02399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06692_ _02329_ _02330_ _02331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_90_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05712_ _01375_ _01337_ _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08500_ _03945_ _03992_ _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09480_ ci_neuron.output_memory\[16\] _04698_ _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05643_ _01247_ _01308_ _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_108_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08431_ _03929_ _03931_ _03932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05703__A1 _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05574_ _01166_ _01199_ _01201_ _01242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08362_ net292 net399 _03871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07313_ _02941_ _02932_ _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08293_ _03796_ net348 _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07244_ _02548_ _02725_ _02874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07175_ _02804_ _02805_ _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06126_ _01779_ _01781_ _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06057_ _01710_ _01711_ _01713_ _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_2_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05008_ internal_ih.byte3\[3\] _00696_ _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06778__I _02415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09816_ _00395_ clknet_leaf_135_sys_clock_i internal_ih.current_instruction\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_129_Left_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06959_ _01850_ _02592_ _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09747_ _00326_ clknet_leaf_33_sys_clock_i ci_neuron.uut_simple_neuron.x2\[28\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09678_ _00265_ clknet_leaf_49_sys_clock_i ci_neuron.uut_simple_neuron.x3\[15\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_83_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08629_ _03900_ _04102_ _04097_ _03892_ _03943_ _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_139_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05170__A2 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_138_Left_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07998__A2 net618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_94_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_125_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08970__I1 internal_ih.byte6\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_93_sys_clock_i_I clknet_4_11_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09427__A2 _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05290_ _00963_ _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_2_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_3_sys_clock_i clknet_4_1_0_sys_clock_i clknet_leaf_3_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_12_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08980_ net373 internal_ih.byte6\[7\] _04257_ _04338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07931_ _03506_ _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07862_ _03446_ _03447_ _03449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06813_ _02447_ _02449_ _02450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09601_ net310 _00555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07793_ net595 _03392_ _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09532_ _04696_ _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06744_ _02223_ _02340_ _02381_ _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_06675_ _02313_ _02274_ _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09463_ net156 _04680_ _04685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05626_ _01289_ _01291_ _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_65_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04846__I _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09394_ ci_neuron.output_val_internal\[3\] _04611_ _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08414_ net647 _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05557_ _01192_ _01224_ _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08345_ net429 net291 _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_22_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05488_ _01157_ _01124_ _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08276_ ci_neuron.uut_simple_neuron.x0\[13\] _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_34_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07227_ _02811_ _02814_ _02856_ _02857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07158_ _02787_ _02788_ _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_113_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06109_ _01713_ _01763_ _01764_ _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_14_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07089_ net38 _02684_ _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06301__I _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_96_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09432__I2 _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_81_sys_clock_i_I clknet_4_14_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06159__A1 ci_neuron.uut_simple_neuron.x2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_85_sys_clock_i clknet_4_14_0_sys_clock_i clknet_leaf_85_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05906__A1 _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06460_ _02103_ _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_87_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05411_ _01048_ _01051_ _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06391_ _01987_ _02034_ _02035_ _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08130_ net614 ci_neuron.uut_simple_neuron.titan_id_0\[21\] _03673_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05342_ _01013_ _01014_ _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_60_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06634__A2 _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05273_ _00946_ _00947_ _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08061_ _03607_ _03612_ _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_60_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07012_ _02641_ _02645_ _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08963_ internal_ih.byte6\[7\] net345 _04327_ _04329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07914_ _03489_ net426 _03492_ _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08894_ net494 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07845_ ci_neuron.uut_simple_neuron.titan_id_2\[4\] net590 _03435_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_07776_ net718 _00110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06570__A1 _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04988_ internal_ih.byte2\[2\] _00686_ _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06727_ _01946_ _01952_ _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09515_ ci_neuron.output_memory\[21\] _04722_ _04729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09446_ _03783_ net84 _00977_ _02139_ _04667_ _04669_ _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_06658_ _02262_ _02297_ _02298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_93_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06589_ _02139_ _02187_ _02229_ _02230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05609_ _01251_ _01275_ _01276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09377_ net180 _04611_ _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08328_ _03840_ _03841_ _03833_ _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_109_sys_clock_i_I clknet_4_8_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08259_ _03781_ _00170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06389__A1 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10221_ _00119_ clknet_leaf_32_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10152_ _00217_ clknet_leaf_40_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[26\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_127_sys_clock_i clknet_4_2_0_sys_clock_i clknet_leaf_127_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_100_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09327__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10083_ _00180_ clknet_leaf_20_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold409 _04272_ net442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_96_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08613__I0 _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09664__D _00251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05960_ net260 _01619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05891_ _01493_ _01551_ _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04911_ internal_ih.byte5\[2\] _00640_ _00641_ internal_ih.byte1\[2\] _00644_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07630_ _02542_ _02562_ _03255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04842_ internal_ih.current_instruction\[0\] internal_ih.current_instruction\[1\]
+ internal_ih.current_instruction\[2\] _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_49_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07561_ _03185_ _03186_ _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_28_sys_clock_i_I clknet_4_7_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06512_ _02077_ _02107_ _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09300_ _04010_ _04546_ _04560_ _00490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07492_ _03047_ _03049_ _03119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_76_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold144_I ci_neuron.output_val_internal\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06443_ _02085_ _02086_ _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_75_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09231_ _04518_ _00463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06374_ _02018_ _02019_ _02020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_fanout12_I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09162_ _04477_ _00435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05325_ _00962_ _00987_ _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08113_ _03657_ net584 _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_142_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08852__I0 internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09093_ net147 _04427_ _04436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05256_ _00907_ _00920_ _00931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08044_ net605 _00091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05187_ _00812_ _00846_ _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05291__A1 _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09995_ _00510_ clknet_leaf_7_sys_clock_i ci_neuron.input_memory\[1\]\[30\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08946_ _04319_ _00377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08877_ _04269_ _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07828_ ci_neuron.uut_simple_neuron.titan_id_2\[0\] net105 _03421_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07759_ net657 ci_neuron.uut_simple_neuron.titan_id_3\[20\] _03364_ _03365_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_6_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09429_ net107 _04655_ _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10204_ _00100_ clknet_leaf_60_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10135_ _00227_ clknet_leaf_55_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10066_ _00193_ clknet_leaf_79_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05110_ _00773_ _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07262__A2 _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06090_ _01744_ _01745_ _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold206 _04158_ net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold217 _00478_ net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold239 _04198_ net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05041_ ci_neuron.address_i\[2\] _00726_ _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold228 ci_neuron.output_memory\[18\] net261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_113_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_16_sys_clock_i_I clknet_4_1_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08800_ _04235_ _00315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06992_ _02625_ _02622_ _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09780_ _00359_ clknet_leaf_0_sys_clock_i internal_ih.byte3\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05943_ _01557_ _01565_ _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08731_ _04173_ _04174_ _04181_ _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08662_ _04124_ _04126_ _04131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07613_ _01850_ _03228_ _03237_ _03238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_96_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05874_ _01528_ _01530_ _01534_ _01535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08593_ ci_neuron.value_i\[21\] _04013_ _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07544_ _03168_ _03169_ _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__08278__A1 _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07475_ _02504_ _03101_ _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06426_ _02026_ _02068_ _02069_ _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_63_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09214_ _04499_ _04509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_101_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08326__I _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06357_ _01960_ _02002_ _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08825__I0 _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09145_ net155 _04469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06288_ _01858_ _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05308_ _00981_ _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_71_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09076_ _04419_ ci_neuron.stream_o\[12\] _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05239_ _00912_ _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08027_ ci_neuron.uut_simple_neuron.titan_id_1\[4\] ci_neuron.uut_simple_neuron.titan_id_0\[4\]
+ _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold762 internal_ih.byte1\[6\] net813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold773 _03570_ net817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold740 ci_neuron.uut_simple_neuron.titan_id_2\[28\] net773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold751 ci_neuron.uut_simple_neuron.titan_id_2\[27\] net784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09250__I0 _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09978_ _00493_ clknet_leaf_70_sys_clock_i ci_neuron.input_memory\[1\]\[13\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_110_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08929_ net517 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09241__I0 _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06755__A1 _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10118_ _00242_ clknet_leaf_43_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_128_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10049_ net121 clknet_leaf_114_sys_clock_i ci_neuron.output_val_internal\[18\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_141_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05590_ _01252_ _01219_ _01256_ _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_34_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07260_ _02326_ _02817_ _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07191_ _02217_ _02237_ _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06211_ _01823_ _01861_ _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06142_ _01700_ _01769_ _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06073_ _01682_ _01684_ _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05246__A1 _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09901_ _00020_ net10 ci_neuron.address_i\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05024_ _00708_ _00709_ _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_41_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold476_I internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09832_ _00411_ clknet_leaf_95_sys_clock_i ci_neuron.output_memory\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09763_ _00342_ clknet_leaf_135_sys_clock_i internal_ih.byte1\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06975_ _02280_ _02441_ _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08714_ internal_ih.spi_rx_byte_i\[1\] internal_ih.spi_rx_byte_i\[0\] internal_ih.spi_rx_byte_i\[2\]
+ _04174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
Xrebuffer21 _02012_ net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05926_ _01576_ _01585_ _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xrebuffer10 _00861_ net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09694_ _00281_ clknet_leaf_9_sys_clock_i ci_neuron.uut_simple_neuron.x3\[31\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05857_ _01412_ _01516_ _01517_ _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08645_ _04116_ net506 _04111_ _04117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08576_ _04056_ _04058_ _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07527_ _03075_ _03117_ _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05788_ _01449_ _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07458_ _03083_ _03084_ _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_81_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06409_ _02047_ _02053_ _02054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07389_ _02676_ _02858_ _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09128_ _04460_ _00418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05237__A1 _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09059_ _04378_ net204 _04404_ _00405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_102_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold581 ci_neuron.uut_simple_neuron.titan_id_1\[21\] net614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold570 ci_neuron.uut_simple_neuron.titan_id_1\[7\] net603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08726__A2 _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold592 _03547_ net625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06737__A1 _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07217__A2 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2_sys_clock_i clknet_4_1_0_sys_clock_i clknet_leaf_2_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_110_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06728__A1 _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06760_ _02376_ _02378_ _02397_ _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06691_ _02286_ _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05711_ _01332_ _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05642_ _01076_ _01234_ _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_108_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08430_ ci_neuron.normalised_stream_write_address\[0\] _03930_ _03927_ _03931_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_47_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05573_ _01166_ _01199_ _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08361_ net292 _03863_ _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_144_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07312_ _02933_ _02940_ _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08292_ ci_neuron.uut_simple_neuron.x0\[15\] _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07243_ _02862_ _02872_ _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_73_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08405__A1 _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07174_ _02731_ _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06125_ _01731_ _01780_ _01728_ _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06056_ _01573_ _01579_ _01712_ _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_78_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05007_ _00699_ _00051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09815_ net280 clknet_leaf_134_sys_clock_i internal_ih.current_instruction\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06958_ _02590_ _02591_ _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09746_ _00325_ clknet_4_4_0_sys_clock_i ci_neuron.uut_simple_neuron.x2\[27\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09677_ _00264_ clknet_4_13_0_sys_clock_i ci_neuron.uut_simple_neuron.x3\[14\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05909_ _01530_ _01534_ _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06889_ _02524_ _00238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_83_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08628_ _03878_ _04081_ _04102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_68_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08559_ _04043_ _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_25_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08644__A1 _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_84_sys_clock_i clknet_4_14_0_sys_clock_i clknet_leaf_84_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07383__A1 _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05697__A1 _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08635__A1 _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09667__D _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer1 _03062_ net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_136_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04952__I _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07610__A2 _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07930_ ci_neuron.uut_simple_neuron.titan_id_2\[17\] ci_neuron.uut_simple_neuron.titan_id_5\[17\]
+ ci_neuron.uut_simple_neuron.titan_id_2\[16\] ci_neuron.uut_simple_neuron.titan_id_5\[16\]
+ _03506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_139_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07861_ _03448_ _00155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07792_ net446 net781 _03391_ _03392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06812_ _02383_ _02448_ _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09600_ ci_neuron.stream_o\[4\] net309 _04795_ _04796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06743_ _02379_ _02380_ _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09531_ _04721_ _04737_ _04741_ _04742_ _00539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__07126__A1 _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06674_ _01899_ _02313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09462_ _04677_ _04683_ _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05625_ _01227_ _01290_ _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_65_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08413_ _03905_ _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09393_ _04603_ _04624_ _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05556_ _01104_ _01223_ _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08535__S _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08344_ _03855_ _00181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05487_ _01156_ _01126_ _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__06101__A2 _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08275_ _03794_ _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07226_ _02803_ _02810_ _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_131_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07157_ _01921_ _02313_ _02714_ _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_120_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05860__A1 _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06108_ _01706_ _01667_ _01710_ _01764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_30_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07088_ net51 _02692_ _02719_ _02720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_30_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06039_ _01374_ _01659_ _01695_ _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07365__A1 _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ _00308_ clknet_leaf_68_sys_clock_i ci_neuron.uut_simple_neuron.x2\[10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_2_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08617__A1 _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05851__A1 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09432__I3 _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_33_sys_clock_i clknet_4_4_0_sys_clock_i clknet_leaf_33_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05410_ _01034_ _01079_ _01080_ _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_126_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06390_ _01993_ _02011_ _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05341_ _00980_ _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05272_ _00944_ _00945_ _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08060_ net561 ci_neuron.uut_simple_neuron.titan_id_0\[9\] _03614_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07011_ _02642_ _02644_ _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08962_ net358 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07913_ net425 ci_neuron.uut_simple_neuron.titan_id_5\[14\] _03492_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08893_ internal_ih.byte3\[1\] net493 _04285_ _04289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07844_ _03431_ _03433_ _03434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07775_ _03376_ _03377_ _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_27_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04987_ _00688_ _00041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06726_ _02362_ _02363_ _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04857__I _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09514_ _04721_ _04723_ _04726_ _04728_ _00536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06657_ _02268_ _02296_ _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07233__I ci_neuron.uut_simple_neuron.x3\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09445_ _04668_ _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05608_ _01257_ _01274_ _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06588_ _02226_ _02228_ _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_75_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09376_ _04610_ _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05539_ _01177_ _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08327_ _03835_ _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08258_ _03777_ _03780_ _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_62_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07209_ _02779_ _02839_ _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_105_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10220_ _00117_ clknet_leaf_4_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[30\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08189_ net772 net566 _03721_ _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_101_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10151_ _00216_ clknet_leaf_40_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05061__A2 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10082_ _00179_ clknet_leaf_22_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08613__I1 _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07329__A1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04910_ _00643_ _00024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05890_ _01500_ _01502_ _01508_ _01495_ _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__09533__I _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04841_ internal_ih.current_instruction\[5\] internal_ih.current_instruction\[4\]
+ internal_ih.current_instruction\[7\] internal_ih.current_instruction\[6\] _00592_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_45_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07560_ _02497_ _03102_ _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_49_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06511_ _02122_ _02153_ _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07491_ _03075_ _03117_ _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05107__A3 _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09230_ _04064_ _03852_ _04514_ _04518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_14_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06442_ _02051_ _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06373_ _01975_ _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09161_ net100 _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05324_ _00966_ _00986_ _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08112_ net583 ci_neuron.uut_simple_neuron.titan_id_0\[18\] _03658_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09092_ net223 _04416_ _04434_ _04435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08043_ _03598_ net604 _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05255_ _00930_ _00201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05186_ _00863_ _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09994_ _00509_ clknet_leaf_7_sys_clock_i ci_neuron.input_memory\[1\]\[29\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08945_ net345 net410 _04317_ _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09443__I _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08876_ net469 _00347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07827_ net409 _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07758_ _03360_ _03362_ _03363_ _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06709_ _02321_ _02347_ _02348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_94_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07689_ net634 _00124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09428_ _04610_ _04655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09359_ _04373_ _04593_ _04594_ _00515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_105_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05806__A1 _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08843__I1 _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07559__A1 _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09548__A2 _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10203_ _00099_ clknet_leaf_58_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10134_ _00226_ clknet_leaf_55_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10065_ _00190_ clknet_leaf_79_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07731__A1 ci_neuron.uut_simple_neuron.titan_id_4\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08834__I1 _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold207 _00286_ net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_25_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold218 ci_neuron.uut_simple_neuron.titan_id_6\[21\] net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05040_ _00722_ _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold229 _04814_ net262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_113_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09003__A4 _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06991_ _02551_ _02624_ _02625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05942_ _01560_ _01590_ _01600_ _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08730_ net256 _04189_ _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05873_ _00739_ _01531_ _01533_ _01474_ _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__09562__I2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08661_ _04124_ _04126_ _04129_ _04130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07612_ _02802_ _03233_ _03236_ _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_89_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08592_ _03848_ _03850_ _04066_ _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_37_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07543_ ci_neuron.uut_simple_neuron.x3\[29\] _03088_ _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07474_ _02812_ _03019_ _03018_ _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_76_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold519_I internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06425_ _02066_ _02067_ _02064_ _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09213_ _03785_ _04489_ _04508_ _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09144_ _04468_ _00426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06356_ ci_neuron.uut_simple_neuron.x3\[8\] _02001_ _02002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__08825__I1 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06287_ _01860_ _01934_ _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_05307_ _00866_ _00976_ _00980_ _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09075_ _04361_ _04419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05238_ _00895_ _00911_ _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xhold730 ci_neuron.uut_simple_neuron.x0\[8\] net763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08026_ net623 _00088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold763 ci_neuron.uut_simple_neuron.titan_id_0\[24\] net796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold741 ci_neuron.input_memory\[1\]\[29\] net809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold752 ci_neuron.uut_simple_neuron.titan_id_2\[26\] net785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05169_ _00846_ _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold785 _00795_ net829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__09250__I1 _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold774 ci_neuron.uut_simple_neuron.x0\[2\] net818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08202__A2 _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09977_ _00492_ clknet_leaf_48_sys_clock_i ci_neuron.input_memory\[1\]\[12\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08928_ net516 internal_ih.byte4\[0\] _04306_ _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08859_ _04269_ _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_54_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_1_sys_clock_i clknet_4_1_0_sys_clock_i clknet_leaf_1_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_118_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10117_ _00241_ clknet_leaf_37_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06755__A2 _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10048_ net135 clknet_leaf_113_sys_clock_i ci_neuron.output_val_internal\[17\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold90 _00519_ net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_141_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06210_ _01858_ _01860_ _01861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_143_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07190_ _02820_ _02794_ _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_27_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06141_ _01754_ _01794_ _01795_ _01796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06072_ _01727_ _01728_ _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_123_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09900_ _00019_ net9 ci_neuron.address_i\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05023_ ci_neuron.instruction_i\[1\] _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_111_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09831_ net141 clknet_leaf_107_sys_clock_i internal_ih.spi_tx_byte_o\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06974_ _02544_ _02565_ _02607_ _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08991__I0 _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09762_ _00341_ clknet_leaf_135_sys_clock_i internal_ih.byte1\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06410__I _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05925_ _01530_ _01584_ _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08713_ _04170_ internal_ih.spi_rx_byte_i\[3\] _04172_ _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
Xrebuffer11 net43 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09693_ _00280_ clknet_leaf_32_sys_clock_i ci_neuron.uut_simple_neuron.x3\[30\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_05856_ _01413_ _01466_ _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xrebuffer22 _00866_ net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_08644_ _04019_ _04113_ _04114_ _04115_ _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_89_sys_clock_i_I clknet_4_11_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05787_ _01124_ _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08575_ _03841_ _04044_ _04057_ _03943_ _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_49_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07526_ _03120_ _03131_ _03151_ _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07457_ ci_neuron.uut_simple_neuron.x3\[27\] _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07388_ _03015_ _03011_ _03016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06408_ _01955_ _02052_ _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_06339_ _01847_ _01984_ _01985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_122_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08423__A2 _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09127_ net248 _04460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05237__A2 _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09058_ net117 _04379_ _04404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08009_ _03569_ _03571_ _03572_ _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold571 _03599_ net604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold560 _03441_ net593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold582 _03673_ net615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_83_sys_clock_i clknet_4_14_0_sys_clock_i clknet_leaf_83_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold593 ci_neuron.stream_o\[25\] net687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06737__A2 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06673__A1 _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06690_ _02285_ _02329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05710_ _01371_ _01373_ _01374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_144_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05641_ _01305_ _01243_ _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08360_ net399 net387 _03869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_53_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07311_ _02936_ _02939_ _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05572_ _01235_ _01239_ _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_67_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04911__B2 internal_ih.byte1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08291_ _03808_ _03809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07242_ _02871_ _02682_ _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_132_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07173_ _02734_ _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06124_ _01682_ _01684_ _01727_ _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_108_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_77_sys_clock_i_I clknet_4_10_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06055_ _01473_ _01577_ _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__04978__A1 internal_ih.byte1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_125_sys_clock_i clknet_4_3_0_sys_clock_i clknet_leaf_125_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05006_ internal_ih.byte3\[2\] _00696_ _00699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09814_ _00393_ clknet_leaf_140_sys_clock_i internal_ih.byte7\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06957_ _02531_ _02537_ _02591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09745_ _00324_ clknet_leaf_32_sys_clock_i ci_neuron.uut_simple_neuron.x2\[26\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06888_ _02521_ _02523_ _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_05908_ _01567_ _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09676_ _00263_ clknet_leaf_50_sys_clock_i ci_neuron.uut_simple_neuron.x3\[13\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05839_ _01498_ _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_90_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_6_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08627_ ci_neuron.value_i\[27\] _04055_ _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08558_ _03821_ _04038_ _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__04902__B2 internal_ih.byte0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04902__A1 internal_ih.byte4\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07509_ _02996_ _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_108_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08489_ ci_neuron.value_i\[6\] _03944_ _03983_ _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_25_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_32_sys_clock_i clknet_4_4_0_sys_clock_i clknet_leaf_32_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_33_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04969__A1 internal_ih.byte1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold390 internal_ih.byte5\[4\] net423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09626__I _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_136_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer2 _01420_ net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_140_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07860_ _03446_ _03447_ _03448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07791_ net780 net787 _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06811_ ci_neuron.uut_simple_neuron.x3\[17\] ci_neuron.uut_simple_neuron.x3\[18\]
+ _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_06742_ _02339_ _02380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09530_ net175 _04727_ _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09461_ _03797_ net74 _01006_ _02228_ _04667_ _04669_ _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_06673_ _01908_ _02273_ _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_65_sys_clock_i_I clknet_4_13_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05624_ ci_neuron.uut_simple_neuron.x2\[19\] ci_neuron.uut_simple_neuron.x2\[20\]
+ _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_80_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09392_ _03730_ net56 _00758_ _01872_ _04622_ _04623_ _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_65_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08412_ _03914_ _00191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05555_ _01096_ _01149_ _01184_ _01223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08343_ _03849_ _03851_ _03854_ _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_46_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08274_ ci_neuron.uut_simple_neuron.x0\[12\] _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_22_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07225_ _02796_ _02853_ _02854_ _02815_ _02819_ _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_117_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05486_ _01130_ _01134_ _01155_ _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_7_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07156_ _02785_ _02786_ _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07087_ _02675_ _02687_ _02719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06107_ _01578_ _01711_ _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_70_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06038_ _01462_ _01660_ _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05376__A1 _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09728_ _00307_ clknet_leaf_49_sys_clock_i ci_neuron.uut_simple_neuron.x2\[9\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_2_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07989_ _03551_ net696 _03555_ _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09181__I _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_134_sys_clock_i_I clknet_4_2_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09659_ net235 net327 _04826_ _04829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_120_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09290__A2 _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_135_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06800__A1 _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_69_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_105_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_138_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05340_ _00811_ net43 _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_78_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09281__A2 _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05271_ _00944_ _00945_ _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_60_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07010_ _02573_ _02643_ _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_53_sys_clock_i_I clknet_4_15_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08961_ internal_ih.byte6\[6\] net357 _04327_ _04328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_87_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07912_ net427 _00132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08892_ _04288_ _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07843_ _03429_ _03432_ _03433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07774_ net717 net610 _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_hold549_I _03349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04986_ internal_ih.byte2\[1\] _00686_ _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06725_ _01929_ _02324_ _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09513_ net166 _04727_ _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06656_ _02271_ _02295_ _02296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09444_ _03935_ _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05607_ _01259_ _01273_ _01274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_94_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05530__A1 _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06587_ _02227_ _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_96_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09375_ _04596_ _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05538_ _01170_ _01196_ _01205_ _01206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_90_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08326_ _03824_ _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05469_ _01042_ _01093_ _01138_ _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08257_ _03778_ _03779_ _03780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07208_ _02835_ _02838_ _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08188_ _03717_ net488 _03720_ _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07139_ _02770_ _00242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07035__A1 _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_122_sys_clock_i_I clknet_4_3_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10150_ _00215_ clknet_leaf_38_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10081_ net545 clknet_leaf_22_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09583__I0 _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_133_Right_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08774__A1 _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10279_ _00572_ clknet_leaf_108_sys_clock_i ci_neuron.stream_o\[21\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04840_ _00591_ internal_ih.got_all_data vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_144_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07490_ _03106_ _03116_ _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06510_ _02124_ _02152_ _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06441_ _02049_ _02085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_62_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_41_sys_clock_i_I clknet_4_7_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06372_ _01972_ _02018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09160_ _04476_ _00434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05323_ _00959_ _00989_ _00995_ _00996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08111_ _03652_ _03654_ _03656_ _03657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09091_ _04356_ _04431_ _04433_ _04411_ _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_32_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05254_ _00926_ _00929_ _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_72_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08042_ net603 ci_neuron.uut_simple_neuron.titan_id_0\[7\] _03599_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_12_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05185_ _00781_ _00838_ _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09557__A3 _04763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08765__A1 _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09993_ _00508_ clknet_leaf_7_sys_clock_i ci_neuron.input_memory\[1\]\[28\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08944_ _04318_ _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09871__D _00062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08875_ internal_ih.byte2\[1\] net468 _04275_ _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07826_ ci_neuron.uut_simple_neuron.titan_id_4\[1\] net408 _03420_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07757_ net532 ci_neuron.uut_simple_neuron.titan_id_3\[19\] _03363_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_04969_ internal_ih.byte1\[2\] _00675_ _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06708_ _02325_ _02328_ _02346_ _02347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_88_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07688_ _03304_ net633 _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_110_sys_clock_i_I clknet_4_8_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06639_ _02230_ _02279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_109_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09427_ _04652_ _04653_ _04654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09358_ _04385_ _04373_ _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_0_sys_clock_i clknet_4_0_0_sys_clock_i clknet_leaf_0_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07256__A1 _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08309_ _03810_ _03825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09289_ _03979_ _04553_ _04554_ _00485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10202_ _00098_ clknet_leaf_58_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10133_ _00225_ clknet_leaf_55_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10064_ _00065_ clknet_leaf_78_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09308__I0 _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09484__A2 _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07495__A1 _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06298__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05402__I _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold208 ci_neuron.stream_enabled net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_4_10_0_sys_clock_i clknet_0_sys_clock_i clknet_4_10_0_sys_clock_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_40_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold219 ci_neuron.uut_simple_neuron.titan_id_6\[27\] net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06233__I _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08747__A1 _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06990_ ci_neuron.uut_simple_neuron.x3\[20\] _02623_ _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__09547__I0 _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05941_ _01563_ _01589_ _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05872_ _01475_ _01532_ _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08660_ net183 internal_ih.spi_tx_byte_o\[7\] _04128_ _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07611_ _03234_ _03235_ _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09562__I3 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08591_ _03849_ _04066_ _03851_ _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07542_ _03166_ _03167_ _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07486__A1 _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07473_ _03099_ _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06424_ _02066_ _02067_ _02064_ _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09212_ _04017_ _04496_ _04508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06355_ ci_neuron.uut_simple_neuron.x3\[9\] _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09143_ net133 _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05306_ _00895_ _00978_ _00979_ _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06286_ _01931_ _01933_ _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_60_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09074_ _04359_ _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05237_ _00750_ _00896_ _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold720 ci_neuron.input_memory\[1\]\[26\] net803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_08025_ net622 ci_neuron.uut_simple_neuron.titan_id_0\[4\] _03584_ _03585_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_102_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05168_ ci_neuron.uut_simple_neuron.x2\[7\] _00846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold764 ci_neuron.uut_simple_neuron.titan_id_0\[27\] net797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold742 ci_neuron.input_memory\[1\]\[2\] net810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold731 ci_neuron.input_memory\[1\]\[0\] net806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold753 ci_neuron.uut_simple_neuron.titan_id_2\[24\] net786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07410__A1 _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_82_sys_clock_i clknet_4_14_0_sys_clock_i clknet_leaf_82_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold786 ci_neuron.uut_simple_neuron.x0\[20\] net830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_12_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold775 ci_neuron.uut_simple_neuron.x0\[30\] net819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_110_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05099_ _00742_ _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09976_ _00491_ clknet_leaf_69_sys_clock_i ci_neuron.input_memory\[1\]\[11\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09454__I _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08927_ _04308_ _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08858_ _04256_ _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07809_ _03391_ _03394_ _03405_ _03406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09879__CLK net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08789_ _04229_ _00310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_130_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05378__B _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07401__A1 _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10116_ _00240_ clknet_leaf_43_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_128_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10047_ net145 clknet_leaf_113_sys_clock_i ci_neuron.output_val_internal\[16\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_42_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold91 ci_neuron.uut_simple_neuron.x0\[10\] net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold80 ci_neuron.output_val_internal\[10\] net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_141_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06140__A1 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06140_ _01792_ _01793_ _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08443__I _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06071_ _01687_ _01688_ _01726_ _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
Xclkbuf_leaf_124_sys_clock_i clknet_4_3_0_sys_clock_i clknet_leaf_124_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05022_ ci_neuron.instruction_i\[0\] _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08599__B _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09274__I _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09830_ _00409_ clknet_leaf_107_sys_clock_i internal_ih.spi_tx_byte_o\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06973_ _02546_ _02564_ _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05508__S _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09761_ _00340_ clknet_leaf_135_sys_clock_i internal_ih.byte1\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05924_ _01577_ _01581_ _01583_ _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08712_ internal_ih.spi_rx_byte_i\[1\] _04143_ _04171_ _04172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xrebuffer12 _02538_ net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08819__S _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09692_ _00279_ clknet_leaf_8_sys_clock_i ci_neuron.uut_simple_neuron.x3\[29\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xrebuffer23 _01966_ net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05855_ _01413_ _01466_ _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08643_ ci_neuron.value_i\[29\] _04013_ _04115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05786_ _01411_ _01442_ _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08574_ _03832_ _04043_ _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07525_ _03123_ _03130_ _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07459__A1 _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07456_ _02937_ _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07387_ _03013_ _02939_ _03014_ _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06407_ _02049_ _02051_ _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_107_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06338_ _01983_ _01984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09126_ _04459_ _00417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06269_ _01909_ _01911_ _01917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_31_sys_clock_i clknet_4_5_0_sys_clock_i clknet_leaf_31_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_20_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09057_ net203 _04381_ _04402_ _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08008_ net613 net776 _03572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold561 ci_neuron.uut_simple_neuron.titan_id_4\[26\] net594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold550 ci_neuron.uut_simple_neuron.titan_id_1\[18\] net583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold572 _03600_ net605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06198__A1 _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold583 _03674_ net616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold594 ci_neuron.stream_o\[30\] net699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09959_ _00474_ clknet_leaf_5_sys_clock_i ci_neuron.uut_simple_neuron.x0\[30\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09184__I _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05173__A2 _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06673__A2 _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07622__A1 _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_15_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05640_ _01244_ _01305_ _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08438__I _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05571_ _01236_ _01237_ _01238_ _01239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_47_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07310_ _02938_ _02863_ _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_86_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08290_ ci_neuron.uut_simple_neuron.x0\[14\] _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07241_ _02870_ _02867_ _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_80_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07172_ _02676_ _02802_ _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07613__A1 _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06123_ _01737_ _01778_ _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_0_sys_clock_i_I clknet_4_0_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06054_ _01706_ _01667_ _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05005_ _00698_ _00050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09813_ _00392_ clknet_leaf_140_sys_clock_i internal_ih.byte7\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06956_ _02534_ _02536_ _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09744_ _00323_ clknet_leaf_32_sys_clock_i ci_neuron.uut_simple_neuron.x2\[25\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_hold746_I ci_neuron.uut_simple_neuron.titan_id_5\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06887_ _02466_ _02468_ _02522_ _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09675_ _00262_ clknet_leaf_50_sys_clock_i ci_neuron.uut_simple_neuron.x3\[12\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_05907_ _01254_ _01566_ _01567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05838_ _01123_ _01499_ _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_90_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08626_ _04100_ _00276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05769_ _01428_ _01429_ _01431_ _01432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08557_ _03822_ _04038_ _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07508_ _03071_ _03134_ _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_135_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08488_ _03945_ _03982_ _03983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_25_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07439_ _02778_ _02980_ net34 _03065_ _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_135_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09109_ _04356_ _04447_ _04449_ _04370_ _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_33_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_107_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_130_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold380 _03317_ net413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold391 _04325_ net424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_125_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_116_Left_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_107_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_125_Left_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xrebuffer3 _01880_ net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07790_ net594 ci_neuron.uut_simple_neuron.titan_id_3\[26\] _03390_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06810_ _02333_ _02389_ _02446_ _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_134_Left_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06741_ _02337_ _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_69_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09552__I _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09460_ ci_neuron.output_memory\[13\] _04675_ _04682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06672_ _02268_ _02296_ _02310_ _02311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08411_ _03910_ _03913_ _03914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05623_ _00747_ _01268_ _01289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09391_ _04606_ _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_129_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05554_ _00742_ _01193_ _01222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08342_ _03852_ _03849_ _03853_ _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__04896__B2 internal_ih.byte0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout28_I net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05485_ _01144_ _01154_ _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08273_ _03793_ _00172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07224_ _02811_ _02814_ _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09426__I2 _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07155_ _02751_ _02757_ _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07086_ _02668_ _02694_ _02717_ _02718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06106_ _01753_ _01761_ _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06037_ _01692_ _01693_ _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_93_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07988_ net785 net695 _03555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06939_ _02515_ _02517_ _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09727_ _00306_ clknet_leaf_68_sys_clock_i ci_neuron.uut_simple_neuron.x2\[8\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_97_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06325__A1 _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09658_ _04828_ _00580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08609_ _04085_ net771 _04086_ _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09589_ _03926_ _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08873__I0 internal_ih.byte2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08625__I0 _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06800__A2 _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08928__I1 internal_ih.byte4\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08553__A2 _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09372__I _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06316__A1 _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08864__I0 net470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05270_ _00751_ _00942_ _00918_ _00909_ _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_71_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08652__S _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08960_ _04311_ _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07911_ _03489_ net426 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08891_ net495 net503 _04285_ _04288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07842_ ci_neuron.uut_simple_neuron.titan_id_2\[3\] ci_neuron.uut_simple_neuron.titan_id_5\[3\]
+ _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07773_ _03372_ _03374_ _03375_ _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04985_ _00687_ _00040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09512_ _04704_ _04727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06724_ _01948_ _02323_ _02362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08827__S _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06655_ _02294_ _02275_ _02295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09443_ _04666_ _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05606_ _01261_ _01272_ _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09374_ _04603_ _04608_ _04609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06586_ ci_neuron.uut_simple_neuron.x3\[13\] _02227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08325_ _03837_ _03838_ _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_145_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05537_ _01172_ _01195_ _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_35_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05468_ _00983_ _01092_ _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08256_ _03755_ _03771_ net195 _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07207_ _02707_ _02836_ _02837_ _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08187_ net487 net801 _03720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07138_ _02764_ _02766_ _02769_ _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_101_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05399_ _01029_ _01027_ _01070_ _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_42_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09457__I _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07069_ _02638_ _02573_ _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_7_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10080_ _00177_ clknet_leaf_22_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09192__I _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06849__A2 _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08472__S _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10278_ _00571_ clknet_leaf_107_sys_clock_i ci_neuron.stream_o\[20\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08526__A2 _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06537__A1 _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06440_ _02054_ _02058_ _02083_ _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_69_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_145_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06371_ _01945_ _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05322_ _00946_ _00988_ _00995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08110_ ci_neuron.uut_simple_neuron.titan_id_1\[17\] ci_neuron.uut_simple_neuron.titan_id_0\[17\]
+ _03656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08462__A1 ci_neuron.value_i\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09090_ _04365_ _04432_ _04433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05253_ _00927_ _00928_ _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08041_ _03596_ _03597_ _03598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_12_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05184_ _00857_ _00860_ net44 _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_81_sys_clock_i clknet_4_14_0_sys_clock_i clknet_leaf_81_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_3_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09992_ _00507_ clknet_leaf_8_sys_clock_i ci_neuron.input_memory\[1\]\[27\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08943_ net357 net431 _04317_ _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08874_ net477 _00346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07825_ net508 _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09190__A2 _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07756_ net532 ci_neuron.uut_simple_neuron.titan_id_3\[19\] _03362_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_04968_ _00677_ _00064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06707_ _02342_ _02345_ _02346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_88_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07687_ net632 ci_neuron.uut_simple_neuron.titan_id_3\[8\] _03305_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09426_ _03770_ net59 _00867_ _01998_ _04644_ _04645_ _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_04899_ _00636_ _00020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09493__A3 _04709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06638_ _02235_ _02238_ _02277_ _02278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06569_ _01863_ _02175_ _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09357_ _04354_ _04592_ _04376_ _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07256__A2 _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09288_ net57 _04549_ _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08308_ _03823_ _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_133_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08239_ _03762_ _03763_ _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_31_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10201_ _00097_ clknet_leaf_58_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10132_ _00224_ clknet_4_15_0_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10063_ net683 clknet_leaf_78_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_0\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07192__A1 _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08819__I0 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05258__A1 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_123_sys_clock_i clknet_4_3_0_sys_clock_i clknet_leaf_123_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_124_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09244__I0 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold209 ci_neuron.uut_simple_neuron.titan_id_6\[5\] net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_141_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05940_ _01599_ _00217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05871_ ci_neuron.uut_simple_neuron.x2\[25\] _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07610_ _02939_ _03170_ _03235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08590_ _02726_ _03941_ _04070_ _00270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07541_ _03084_ ci_neuron.uut_simple_neuron.x3\[28\] _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07472_ _03080_ _03098_ _03099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06423_ _02016_ _02022_ _02067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_57_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09211_ _04010_ _04503_ _04507_ _00454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06354_ _01959_ _01965_ _01999_ _02000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_84_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09142_ _04467_ _00425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05305_ _00910_ _00977_ _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09483__I0 _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06285_ _01878_ _01932_ _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xclkbuf_leaf_30_sys_clock_i clknet_4_4_0_sys_clock_i clknet_leaf_30_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09073_ _04361_ _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05236_ _00895_ _00911_ _00912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold721 _01184_ net754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09235__I0 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold710 _03689_ net743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08024_ _03580_ _03582_ _03583_ _03584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_13_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold754 ci_neuron.uut_simple_neuron.titan_id_3\[25\] net787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05167_ _00845_ _00225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold732 _02387_ net765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_hold776_I ci_neuron.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold743 net826 net776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold776 ci_neuron.uut_simple_neuron.x3\[0\] net820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold765 _03703_ net798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold787 ci_neuron.uut_simple_neuron.titan_id_6\[26\] net831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_05098_ _00763_ _00771_ _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09975_ _00490_ clknet_leaf_70_sys_clock_i ci_neuron.input_memory\[1\]\[10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08926_ net410 net492 _04306_ _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08857_ _04268_ _00339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07808_ ci_neuron.uut_simple_neuron.titan_id_4\[26\] ci_neuron.uut_simple_neuron.titan_id_3\[26\]
+ _03405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08788_ _04023_ _00971_ _04225_ _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07739_ ci_neuron.uut_simple_neuron.titan_id_4\[17\] ci_neuron.uut_simple_neuron.titan_id_3\[17\]
+ _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09409_ _04627_ _04635_ _04637_ _04638_ _00521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_118_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06988__A1 _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_49_sys_clock_i clknet_4_13_0_sys_clock_i clknet_leaf_49_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09226__I0 _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10115_ _00239_ clknet_leaf_43_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_54_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10046_ net110 clknet_leaf_113_sys_clock_i ci_neuron.output_val_internal\[15\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold92 internal_ih.spi_tx_byte_o\[0\] net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold70 ci_neuron.output_val_internal\[11\] net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold81 _00526_ net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04923__B1 _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06979__A1 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06070_ _01687_ _01688_ _01726_ _01727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09217__I0 _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05021_ _00707_ _00065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09393__A2 _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06972_ _02599_ _02605_ _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_77_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09760_ _00339_ clknet_leaf_131_sys_clock_i internal_ih.byte1\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05923_ _00738_ _01582_ _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09691_ _00278_ clknet_leaf_31_sys_clock_i ci_neuron.uut_simple_neuron.x3\[28\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08711_ internal_ih.spi_rx_byte_i\[7\] internal_ih.spi_rx_byte_i\[6\] internal_ih.spi_rx_byte_i\[5\]
+ internal_ih.spi_rx_byte_i\[4\] _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_83_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08642_ _03900_ _03912_ _04102_ _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xrebuffer13 _02518_ net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_117_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer24 net164 net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_05854_ _01513_ _01514_ _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05785_ _01447_ _00214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08573_ ci_neuron.value_i\[18\] _04055_ _04056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07524_ _03148_ _03149_ _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07459__A2 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07455_ _02859_ _03010_ _03081_ _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06406_ _01964_ _02050_ _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07386_ _02933_ _02940_ _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06337_ _01830_ _01877_ _01982_ _01983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09125_ net160 _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06268_ _01912_ _01914_ _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09208__I0 _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09056_ _04382_ _04399_ _04401_ _04354_ _04402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_32_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05642__A1 _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05219_ _00895_ _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08007_ net613 net776 _03571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold562 _03390_ net595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_06199_ _01836_ net751 _01846_ _01850_ _00164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold551 _03658_ net584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold540 ci_neuron.uut_simple_neuron.titan_id_1\[5\] net573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06198__A2 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold584 ci_neuron.uut_simple_neuron.x0\[18\] net617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold573 ci_neuron.uut_simple_neuron.titan_id_1\[3\] net606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold595 ci_neuron.stream_o\[2\] net700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09958_ _00473_ clknet_leaf_5_sys_clock_i ci_neuron.uut_simple_neuron.x0\[29\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08909_ net490 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07147__A1 _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09889_ _00050_ net18 ci_neuron.value_i\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_128_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_56_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09375__I _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10029_ net95 clknet_leaf_7_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05570_ _01169_ _01197_ _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_47_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07240_ _02797_ _02869_ _02870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_80_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__04982__I _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07171_ _02799_ _02801_ _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05872__A1 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06122_ _01594_ _01777_ _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09869__CLK net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06053_ _01473_ _01577_ _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05004_ internal_ih.byte3\[1\] _00696_ _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09812_ _00391_ clknet_leaf_142_sys_clock_i internal_ih.byte7\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_90_sys_clock_i_I clknet_4_11_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07129__A1 _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06955_ _02589_ _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09743_ _00322_ clknet_leaf_32_sys_clock_i ci_neuron.uut_simple_neuron.x2\[24\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06886_ _02408_ _02406_ _02463_ _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09674_ _00261_ clknet_leaf_50_sys_clock_i ci_neuron.uut_simple_neuron.x3\[11\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05906_ _01179_ _01565_ _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05837_ _01496_ _01305_ _01498_ _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08625_ _04099_ _03083_ _04086_ _04100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_96_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08556_ _04041_ _00265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07507_ _03073_ _03133_ _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05768_ _01344_ _01430_ _01431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08629__B2 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05699_ _01341_ _01346_ _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08487_ _03753_ _03976_ _03982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07438_ _03059_ _03063_ _03064_ _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_135_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07369_ _02924_ _02949_ _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09108_ _04365_ _04448_ _04449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_49_sys_clock_i_I clknet_4_13_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09039_ _04358_ ci_neuron.stream_o\[9\] _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold381 ci_neuron.uut_simple_neuron.titan_id_5\[21\] net414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold370 internal_ih.byte5\[1\] net403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold392 ci_neuron.uut_simple_neuron.titan_id_2\[14\] net425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06040__A1 _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09380__I2 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07540__A1 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09293__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer4 net36 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_118_sys_clock_i_I clknet_4_6_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10191__D _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06740_ _02342_ _02345_ _02377_ _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_69_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06671_ _02271_ _02295_ _02310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_78_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05622_ _00750_ _01287_ _01270_ _01263_ _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_08410_ _03907_ _03911_ net418 _03906_ _03913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_74_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09390_ _04604_ _04622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09659__I0 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05553_ _01218_ _01220_ _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08341_ _03844_ _03846_ _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05484_ _01153_ _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08272_ _03789_ _03792_ _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_62_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_22_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07223_ _02811_ _02814_ _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_117_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08882__I1 net470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09426__I3 _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07154_ _02754_ _02756_ _02785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07598__A1 _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09587__A2 _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07085_ _02671_ _02693_ _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold591_I ci_neuron.uut_simple_neuron.titan_id_5\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06105_ _01714_ _01760_ _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06270__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06036_ _01568_ _01677_ _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05048__I net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07987_ ci_neuron.uut_simple_neuron.titan_id_2\[27\] net618 _03554_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06938_ _02569_ _02572_ _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09726_ _00305_ clknet_leaf_66_sys_clock_i ci_neuron.uut_simple_neuron.x2\[7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_9_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09511__A2 _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06869_ _02497_ _02504_ _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08570__I0 _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09657_ net223 net196 _04826_ _04828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_37_sys_clock_i_I clknet_4_5_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08608_ _03939_ _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09588_ _00710_ _00713_ _00725_ _04788_ _00550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_120_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08539_ ci_neuron.value_i\[13\] _04025_ _04026_ _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_41_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09027__A1 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08625__I1 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06013__A1 _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_109_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_106_sys_clock_i_I clknet_4_8_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08732__I _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09569__A2 _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_80_sys_clock_i clknet_4_14_0_sys_clock_i clknet_leaf_80_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_12_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07910_ net425 ci_neuron.uut_simple_neuron.titan_id_5\[14\] _03490_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08890_ _04287_ _00353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07841_ net608 net735 _03431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07772_ net640 ci_neuron.uut_simple_neuron.titan_id_3\[22\] _03375_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06723_ _02319_ _02348_ _02360_ _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_04984_ internal_ih.byte2\[0\] _00686_ _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09511_ _04724_ _04725_ _04726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06654_ _02278_ _02293_ _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_78_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ _03930_ _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06585_ net500 _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05605_ _01262_ _01271_ _01272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09373_ _03725_ net86 _00736_ _02898_ _04605_ _04607_ _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_05536_ _01204_ _00208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08324_ _03835_ net393 _03838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05818__A1 _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05467_ _01083_ _01135_ _01136_ _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__10096__D _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08255_ net195 net578 _03761_ _03764_ _03765_ _03778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_07206_ _02709_ _02760_ _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05398_ _01065_ _01069_ _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08186_ _03719_ _00086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07137_ _02767_ _02768_ _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_99_sys_clock_i clknet_4_10_0_sys_clock_i clknet_leaf_99_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_113_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07068_ _02576_ _02641_ _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06019_ _01657_ _01676_ _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_25_sys_clock_i_I clknet_4_6_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09709_ net149 clknet_leaf_105_sys_clock_i internal_ih.spi_rx_byte_i\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05809__A1 _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_sys_clock_i sys_clock_i clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_52_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_122_sys_clock_i clknet_4_3_0_sys_clock_i clknet_leaf_122_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_133_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10277_ _00570_ clknet_leaf_108_sys_clock_i ci_neuron.stream_o\[19\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07734__A1 _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06537__A2 _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08782__I0 _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_144_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06370_ _02015_ _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05321_ _00953_ _00956_ _00991_ _00951_ _00994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_32_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05252_ _00851_ _00875_ _00882_ _00902_ _00877_ _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_08040_ _03593_ _03594_ _03597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_12_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09558__I _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06225__A1 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05183_ ci_neuron.uut_simple_neuron.x2\[7\] ci_neuron.uut_simple_neuron.x2\[8\] _00861_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_4_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09991_ _00506_ clknet_leaf_33_sys_clock_i ci_neuron.input_memory\[1\]\[26\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08942_ _04311_ _04317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_86_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08873_ internal_ih.byte2\[0\] net476 _04275_ _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07824_ net507 ci_neuron.uut_simple_neuron.titan_id_3\[31\] _03418_ _03419_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07755_ net533 _00105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04967_ internal_ih.byte1\[1\] _00675_ _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06706_ _02344_ _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07686_ _03302_ _03303_ _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_88_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold721_I _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06637_ _02225_ _02276_ _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04898_ internal_ih.byte4\[5\] _00633_ _00634_ internal_ih.byte0\[5\] _00636_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09425_ _04602_ _04652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06568_ _02203_ _02205_ _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09356_ _04145_ _04179_ _04385_ _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06499_ ci_neuron.uut_simple_neuron.x3\[12\] _02142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05519_ _01186_ _01187_ _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xclkbuf_leaf_48_sys_clock_i clknet_4_6_0_sys_clock_i clknet_leaf_48_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09287_ _04543_ _04553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08307_ net406 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_144_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08238_ _03752_ ci_neuron.uut_simple_neuron.x0\[7\] _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10200_ _00126_ clknet_leaf_58_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_5\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08169_ net680 ci_neuron.uut_simple_neuron.titan_id_0\[28\] _03705_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10131_ _00223_ clknet_leaf_63_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10062_ net245 clknet_leaf_123_sys_clock_i ci_neuron.output_val_internal\[31\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_8_sys_clock_i_I clknet_4_4_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08819__I1 _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09244__I1 _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09547__I2 _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05870_ ci_neuron.uut_simple_neuron.x2\[24\] ci_neuron.uut_simple_neuron.x2\[25\]
+ _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07540_ _03083_ _03088_ _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04941__A1 internal_ih.byte6\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07471_ _03093_ _03097_ _03098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_17_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06422_ _01981_ _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09210_ _04005_ _04496_ _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06353_ _01960_ _01998_ _01999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09141_ net265 _04467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05304_ _00910_ _00977_ _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_71_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09072_ _04370_ _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06284_ ci_neuron.uut_simple_neuron.x3\[6\] ci_neuron.uut_simple_neuron.x3\[7\] _01932_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_71_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08023_ net606 ci_neuron.uut_simple_neuron.titan_id_0\[3\] _03583_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_10_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05235_ net759 _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold711 ci_neuron.input_memory\[1\]\[15\] net793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_53_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold700 internal_ih.current_instruction\[1\] net733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05166_ _00830_ _00831_ _00844_ _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xhold722 _01052_ net755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold744 ci_neuron.uut_simple_neuron.titan_id_0\[20\] net777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold733 ci_neuron.uut_simple_neuron.titan_id_3\[0\] net807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold755 ci_neuron.uut_simple_neuron.titan_id_0\[26\] net788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_12_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold777 ci_neuron.input_memory\[1\]\[12\] net821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold766 ci_neuron.uut_simple_neuron.titan_id_1\[29\] net799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05097_ _00736_ _00774_ _00772_ _00775_ _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_09974_ _00489_ clknet_leaf_74_sys_clock_i ci_neuron.input_memory\[1\]\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08925_ _04307_ _00368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05056__I _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08856_ net468 net501 _04264_ _04268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07807_ _03390_ _03403_ _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05999_ _01655_ _01656_ _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08787_ _04228_ _00309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07738_ net581 _03346_ _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07669_ net631 _00121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06685__A1 _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05488__A2 _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09408_ net177 _04633_ _04638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09339_ _04582_ _00507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_117_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09198__I _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08426__A2 _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10114_ _00238_ clknet_leaf_44_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_112_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10132__CLK clknet_4_15_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10045_ net116 clknet_leaf_113_sys_clock_i ci_neuron.output_val_internal\[14\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold60 ci_neuron.input_memory\[1\]\[28\] net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold71 _00527_ net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold82 ci_neuron.output_val_internal\[14\] net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_89_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold93 _04144_ net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_141_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04923__B2 internal_ih.byte1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05020_ net32 _00706_ _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06971_ _02602_ _02604_ _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05922_ _01533_ _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09690_ _00277_ clknet_leaf_25_sys_clock_i ci_neuron.uut_simple_neuron.x3\[27\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08710_ net227 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05853_ _01456_ _01488_ _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08641_ _03915_ _04107_ _04113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xrebuffer14 net46 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer25 _02145_ net274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_05784_ _01444_ _01446_ _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08572_ _03950_ _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07523_ _03071_ _03134_ _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_88_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07454_ _03007_ _03009_ _03081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_hold517_I ci_neuron.uut_simple_neuron.x2\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06405_ ci_neuron.uut_simple_neuron.x3\[9\] ci_neuron.uut_simple_neuron.x3\[10\]
+ _02050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_17_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07385_ _03012_ _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_106_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06336_ _01835_ _01952_ _01982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09124_ _04458_ _00416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06267_ _01915_ _00167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09055_ _04389_ _04400_ _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05218_ ci_neuron.uut_simple_neuron.x2\[9\] _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold530 _03613_ net563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08006_ net817 _00148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06198_ _01847_ _01848_ _01849_ _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_102_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold552 _03659_ net585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold541 _03589_ net574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold563 net69 net683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07395__A2 _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06198__A3 _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05149_ _00828_ _00224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold596 ci_neuron.uut_simple_neuron.titan_id_3\[5\] net629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold585 ci_neuron.uut_simple_neuron.titan_id_5\[27\] net618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold574 _03581_ net607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09957_ _00472_ clknet_leaf_6_sys_clock_i ci_neuron.uut_simple_neuron.x0\[28\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08908_ internal_ih.byte3\[7\] net489 _04296_ _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09392__I0 _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09888_ _00049_ net18 ci_neuron.value_i\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08839_ net501 _04146_ _04258_ _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05881__A2 _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput4 net4 spi_poci_o vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_31_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09391__I _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10028_ net93 clknet_leaf_5_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[30\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07170_ _02730_ _02800_ _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09063__A2 ci_neuron.stream_o\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06121_ _01740_ _01776_ _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06052_ _01707_ _01708_ _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05624__A2 ci_neuron.uut_simple_neuron.x2\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08470__I _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05003_ _00697_ _00049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07377__A2 _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09811_ _00390_ clknet_leaf_141_sys_clock_i internal_ih.byte7\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09742_ _00321_ clknet_leaf_31_sys_clock_i ci_neuron.uut_simple_neuron.x2\[23\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_06954_ _02576_ _02588_ _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06885_ net46 _02520_ _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_118_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09673_ _00260_ clknet_leaf_51_sys_clock_i ci_neuron.uut_simple_neuron.x3\[10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05905_ _01419_ _01420_ _01525_ _01564_ _01429_ _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_05836_ _01304_ _01355_ _01497_ _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_90_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08624_ _04055_ _04096_ _04097_ _04098_ _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05767_ _01328_ _01382_ _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08555_ _04040_ net765 _04028_ _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07506_ _03118_ _03132_ _03133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05560__A1 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05698_ _01218_ _01325_ _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08486_ _03957_ _03979_ _03981_ _00255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07437_ _02983_ _03062_ _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_135_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07368_ _02994_ _02971_ _02995_ _02996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_134_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06165__I ci_neuron.uut_simple_neuron.x3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06319_ _01965_ _01903_ _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09107_ ci_neuron.output_val_internal\[31\] ci_neuron.output_val_internal\[23\] ci_neuron.output_val_internal\[15\]
+ ci_neuron.output_val_internal\[7\] _04366_ _04367_ _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_115_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07299_ ci_neuron.uut_simple_neuron.x3\[23\] _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09038_ _04360_ _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold360 ci_neuron.uut_simple_neuron.x0\[19\] net393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold371 spi_interface_cvonk.state\[0\] net404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold393 _03490_ net426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08565__A1 _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold382 _03523_ net415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09380__I3 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer5 _02678_ net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_7_0_sys_clock_i clknet_0_sys_clock_i clknet_4_7_0_sys_clock_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_20_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_39_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_69_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06670_ _02256_ _02299_ _02309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05621_ _01226_ ci_neuron.uut_simple_neuron.x2\[19\] _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05552_ _00886_ _01207_ _01219_ _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_73_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08340_ _03836_ _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_50_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05483_ _01133_ _01152_ _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_80_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08271_ _03790_ _03791_ _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_11_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07222_ _02821_ _02831_ _02851_ _02852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07153_ _02716_ _02782_ _02783_ _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_116_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06104_ _01756_ _01759_ _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_98_sys_clock_i clknet_4_10_0_sys_clock_i clknet_leaf_98_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07084_ _02712_ _02715_ _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06035_ _01657_ _01676_ _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08547__A1 _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07986_ _03553_ _00145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06937_ _02570_ _02514_ _02571_ _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09725_ _00304_ clknet_leaf_66_sys_clock_i ci_neuron.uut_simple_neuron.x2\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09347__I0 _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09656_ _04827_ _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06868_ _02380_ _02503_ _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__05064__I _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08570__I1 _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08607_ _04019_ _04082_ _04083_ _04084_ _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XANTENNA__05533__A1 _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06799_ _02135_ _02394_ _02435_ _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_05819_ _01479_ _01480_ _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09587_ _00710_ _00713_ net138 _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08538_ _03943_ _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_41_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08469_ _03963_ _03964_ _03966_ _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA_clkbuf_4_8_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_121_sys_clock_i clknet_4_3_0_sys_clock_i clknet_leaf_121_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_135_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06261__A2 _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold190 ci_neuron.stream_o\[29\] net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__09338__I0 _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08777__A1 _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06252__A2 _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07840_ net609 _00152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07771_ net640 ci_neuron.uut_simple_neuron.titan_id_3\[22\] _03374_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_75_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09329__I0 _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06722_ _02321_ _02347_ _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09510_ _03848_ ci_neuron.input_memory\[1\]\[20\] ci_neuron.uut_simple_neuron.x2\[20\]
+ _02620_ _04716_ _04717_ _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XPHY_EDGE_ROW_56_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_04983_ _00685_ _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07504__A2 _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06653_ _02289_ _02292_ _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09441_ ci_neuron.output_memory\[11\] _04650_ _04665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06584_ _02086_ _02189_ _02224_ _02225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05604_ _01263_ _01270_ _01271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout33_I ci_neuron.uut_simple_neuron.x2\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09372_ _04606_ _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05535_ _01200_ _01203_ _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08323_ _03835_ _03836_ _03837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_47_sys_clock_i clknet_4_6_0_sys_clock_i clknet_leaf_47_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_75_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05466_ _01090_ _01094_ _01136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08254_ net578 _03776_ _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__08923__I _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07205_ _02709_ _02760_ _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05397_ _01066_ _01023_ _01068_ _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_65_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08185_ _03717_ net488 _03719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07136_ _02639_ _02637_ _02765_ _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_132_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08768__A1 _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07067_ _02648_ _02699_ _02700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_3_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06018_ _01661_ _01675_ _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05059__I _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09568__I0 _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09193__A1 _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_74_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09708_ net202 clknet_leaf_105_sys_clock_i internal_ih.spi_rx_byte_i\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07969_ ci_neuron.uut_simple_neuron.titan_id_2\[23\] net497 ci_neuron.uut_simple_neuron.titan_id_2\[22\]
+ net458 _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_97_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09496__A2 _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09639_ net471 ci_neuron.output_memory\[21\] _04816_ _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08833__I _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06234__A2 _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10276_ _00569_ clknet_leaf_107_sys_clock_i ci_neuron.stream_o\[18\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08782__I1 _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05320_ _00960_ _00990_ _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05251_ _00882_ _00902_ _00927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_83_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__04859__I0 internal_ih.byte4\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05182_ _00859_ _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06225__A2 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09990_ _00505_ clknet_leaf_31_sys_clock_i ci_neuron.input_memory\[1\]\[25\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08941_ net422 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08872_ net479 _00345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold282_I ci_neuron.output_memory\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07823_ _03414_ _03416_ _03417_ _03418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07094__I _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07754_ net532 ci_neuron.uut_simple_neuron.titan_id_3\[19\] _03360_ _03361_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_04966_ _00676_ _00063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06705_ _02085_ _02343_ _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_07685_ _03299_ _03300_ _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_88_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06636_ _02136_ _02233_ _02276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04897_ _00635_ _00019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09424_ ci_neuron.output_memory\[8\] _04650_ _04651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06567_ _02208_ _00232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09355_ _04591_ _00514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06498_ _02089_ _02095_ _02140_ _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05518_ _01096_ ci_neuron.uut_simple_neuron.x2\[16\] ci_neuron.uut_simple_neuron.x2\[17\]
+ _01187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_63_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09286_ _03974_ _04544_ _04552_ _00484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08306_ _03821_ _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05449_ _01119_ _01071_ _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_90_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08237_ _03741_ _03752_ _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08168_ _03692_ _03700_ net798 _03704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07119_ _02749_ _02750_ _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08099_ net586 net546 _03647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10130_ _00200_ clknet_leaf_63_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_3\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10061_ net259 clknet_leaf_123_sys_clock_i ci_neuron.output_val_internal\[30\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05727__A1 _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_98_sys_clock_i_I clknet_4_10_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07404__A1 _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07955__A2 ci_neuron.uut_simple_neuron.titan_id_5\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09547__I3 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10259_ _00552_ clknet_leaf_95_sys_clock_i ci_neuron.stream_o\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07470_ _02725_ _03096_ _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06421_ _02065_ _00229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06352_ _01964_ _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09140_ _04466_ _00424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_57_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06283_ _01874_ _01904_ _01930_ _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05303_ ci_neuron.uut_simple_neuron.x2\[11\] _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09483__I2 _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09071_ _04377_ _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08022_ net606 ci_neuron.uut_simple_neuron.titan_id_0\[3\] _03582_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_141_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05234_ ci_neuron.uut_simple_neuron.x2\[10\] _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold712 ci_neuron.input_memory\[1\]\[18\] net794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold701 _00476_ net734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05165_ _00834_ _00843_ _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold734 _00753_ net767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold723 ci_neuron.uut_simple_neuron.x3\[28\] net756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold745 _03669_ net778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout5 net8 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05096_ _00777_ _00200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold767 ci_neuron.uut_simple_neuron.titan_id_2\[15\] net800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09973_ _00488_ clknet_leaf_67_sys_clock_i ci_neuron.input_memory\[1\]\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold778 ci_neuron.uut_simple_neuron.x0\[9\] net822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold756 ci_neuron.uut_simple_neuron.titan_id_2\[25\] net789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08924_ net431 net482 _04306_ _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08855_ _04267_ _00338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07806_ _03397_ _03399_ _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08786_ _04017_ net752 _04225_ _04228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07737_ _03342_ _03343_ _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05998_ _01527_ _01626_ _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04949_ internal_ih.byte0\[1\] _00665_ _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_138_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07668_ _03287_ net630 _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06685__A2 _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07599_ _02604_ _02630_ _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06619_ _01836_ _02212_ _02259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09407_ _04630_ _04636_ _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09338_ _04104_ net72 _04578_ _04582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09479__I _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07634__A1 _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09269_ _04139_ _04535_ net300 _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09387__A1 ci_neuron.output_val_internal\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_86_sys_clock_i_I clknet_4_14_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10113_ _00237_ clknet_leaf_43_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_112_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10044_ net157 clknet_leaf_116_sys_clock_i ci_neuron.output_val_internal\[13\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold50 _00518_ net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold61 net807 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold83 _00530_ net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold72 ci_neuron.uut_simple_neuron.titan_id_5\[0\] net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold94 ci_neuron.output_val_internal\[12\] net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_141_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07625__A1 _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08976__I1 internal_ih.byte6\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06970_ _02125_ _02127_ _02603_ _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_05921_ _01574_ _01578_ _01580_ _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05852_ _01460_ _01487_ _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08640_ _04112_ _00278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer15 _02641_ net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer26 _02288_ net318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_05783_ _01400_ _01404_ _01445_ _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_85_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08571_ _04054_ _00267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07522_ _03073_ _03147_ _03148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07453_ _03011_ _03015_ _03079_ _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06404_ _01961_ _02002_ _02048_ _02049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_17_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07384_ _02936_ _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09123_ net242 _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07616__A1 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06335_ _01976_ _01978_ _01981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_33_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06266_ _01912_ _01914_ _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09054_ ci_neuron.output_val_internal\[26\] ci_neuron.output_val_internal\[18\] ci_neuron.output_val_internal\[10\]
+ ci_neuron.output_val_internal\[2\] _04390_ _04391_ _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_44_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05217_ _00869_ _00893_ _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold520 ci_neuron.uut_simple_neuron.titan_id_2\[31\] net553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08005_ net613 net776 _03569_ _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
Xhold542 ci_neuron.uut_simple_neuron.titan_id_4\[21\] net575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_06197_ _01837_ _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold553 ci_neuron.uut_simple_neuron.titan_id_1\[15\] net586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold531 ci_neuron.uut_simple_neuron.titan_id_2\[8\] net564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05148_ _00806_ _00827_ _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold597 _03288_ net630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold575 ci_neuron.uut_simple_neuron.titan_id_2\[3\] net608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold564 ci_neuron.uut_simple_neuron.titan_id_0\[0\] net686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold586 _03554_ net619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_110_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05067__I _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05079_ _00759_ _00761_ _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09956_ _00471_ clknet_leaf_6_sys_clock_i ci_neuron.uut_simple_neuron.x0\[27\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08907_ net467 _00360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09887_ _00048_ net17 ci_neuron.value_i\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08838_ _04257_ _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_142_Right_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08769_ _03974_ _04209_ _04217_ _00302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_74_sys_clock_i_I clknet_4_12_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05094__A1 _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10027_ net72 clknet_leaf_7_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06897__A2 _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_143_sys_clock_i_I clknet_4_0_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_97_sys_clock_i clknet_4_10_0_sys_clock_i clknet_leaf_97_sys_clock_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06120_ _01743_ _01775_ _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06051_ _01618_ _01620_ _01671_ _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_124_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05002_ internal_ih.byte3\[0\] _00696_ _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09810_ _00389_ clknet_leaf_137_sys_clock_i internal_ih.byte7\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06953_ _02587_ _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09741_ _00320_ clknet_leaf_31_sys_clock_i ci_neuron.uut_simple_neuron.x2\[22\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05904_ _01427_ _01525_ _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06884_ _02464_ _02462_ _02519_ _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09672_ _00259_ clknet_leaf_69_sys_clock_i ci_neuron.uut_simple_neuron.x3\[9\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05835_ _01400_ _01444_ _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
X_08623_ ci_neuron.value_i\[26\] _03965_ _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05766_ _01423_ _01419_ _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08554_ _03996_ _04037_ _04038_ _04039_ _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_07505_ _03120_ _03131_ _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05560__A2 _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05697_ _01254_ _01325_ _01360_ _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08485_ net769 _03980_ _03981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07436_ _02991_ _02988_ _03063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10122__CLK clknet_4_5_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_120_sys_clock_i clknet_4_3_0_sys_clock_i clknet_leaf_120_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07367_ _02922_ _02961_ _02995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_116_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06318_ _01960_ _01964_ _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_98_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09106_ _04417_ ci_neuron.stream_o\[7\] ci_neuron.stream_o\[23\] _04418_ _04446_
+ _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_32_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07298_ _02731_ _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09037_ _04359_ _04384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06249_ _01830_ _01881_ _01897_ _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_102_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold361 internal_ih.expected_byte_count\[0\] net394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold350 ci_neuron.uut_simple_neuron.titan_id_6\[2\] net383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold394 _03491_ net427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold383 _03524_ net416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold372 _00477_ net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_leaf_62_sys_clock_i_I clknet_4_14_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09939_ _00454_ clknet_leaf_73_sys_clock_i ci_neuron.uut_simple_neuron.x0\[10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08836__I _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09373__S0 _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_139_sys_clock_i clknet_4_0_0_sys_clock_i clknet_leaf_139_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_126_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer6 _02772_ net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_140_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_131_sys_clock_i_I clknet_4_2_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05620_ _01261_ _01272_ _01285_ _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07650__I _03274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05551_ _01105_ _01151_ _01192_ _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05482_ _01148_ _01151_ _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08270_ _03782_ _03784_ _03786_ _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07221_ _02794_ _02820_ _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08619__I0 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07152_ _02718_ _02759_ _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06103_ _01669_ _01757_ _01758_ _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07083_ _01835_ _01871_ _02714_ _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_124_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06034_ _01689_ _01690_ _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07985_ _03551_ net696 _03553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06936_ _02474_ _02513_ _02571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05345__I _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09724_ _00303_ clknet_leaf_66_sys_clock_i ci_neuron.uut_simple_neuron.x2\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06867_ _02500_ _02502_ _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_2_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09655_ net152 net198 _04826_ _04827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_145_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05818_ _01433_ _01291_ _01380_ _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08606_ ci_neuron.value_i\[23\] _04013_ _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06798_ _02096_ _02279_ _02435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09586_ _04787_ _00549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_120_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05749_ _01255_ _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08537_ _03797_ _03798_ _04015_ _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_41_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08468_ ci_neuron.value_i\[3\] _03965_ _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08483__A1 ci_neuron.value_i\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07419_ _01867_ _01936_ _03045_ _03046_ _03047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_108_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_50_sys_clock_i_I clknet_4_13_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08399_ ci_neuron.uut_simple_neuron.x0\[28\] _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09283__I0 _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold180 ci_neuron.output_val_internal\[1\] net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07735__I net694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold191 _04435_ net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_137_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07277__A2 _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05288__A1 _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09397__I _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06788__A1 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07770_ net641 _00109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04982_ _00599_ _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06721_ _02315_ _02316_ _02317_ _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_3_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09440_ _04649_ _04661_ _04663_ _04664_ _00526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06652_ _02291_ _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06583_ _02222_ _02223_ _02224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05603_ _00741_ _01265_ _01269_ _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_75_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09371_ _03935_ _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05534_ _01201_ _01202_ _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08322_ net393 _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout26_I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08253_ net124 _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07204_ _02781_ _02834_ _02835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_117_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05465_ _01090_ _01094_ _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05396_ _01067_ _01024_ _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08184_ net487 ci_neuron.uut_simple_neuron.titan_id_0\[30\] _03718_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07135_ _02700_ _02705_ _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_hold694_I _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07066_ _02649_ _02698_ _02699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06017_ _01674_ _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_7_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09193__A2 _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05203__A1 _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07968_ _03531_ _03536_ _03538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06919_ _02445_ _02501_ _02553_ _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09707_ net240 clknet_leaf_106_sys_clock_i internal_ih.spi_rx_byte_i\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07899_ _03477_ _03479_ _03480_ _03481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_69_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06703__A1 _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09638_ net324 _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_104_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09569_ _04768_ _04774_ _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08456__A1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09256__I0 _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10275_ _00568_ clknet_leaf_109_sys_clock_i ci_neuron.stream_o\[17\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05250_ _00922_ _00925_ _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_72_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04859__I1 internal_ih.byte3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05181_ _00858_ _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_12_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_90_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08940_ net421 internal_ih.byte4\[5\] _04312_ _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08871_ internal_ih.byte1\[7\] net478 _04275_ _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07822_ ci_neuron.uut_simple_neuron.titan_id_4\[30\] ci_neuron.uut_simple_neuron.titan_id_3\[30\]
+ _03417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07753_ _03350_ _03355_ _03356_ _03358_ _03359_ _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_04965_ internal_ih.byte1\[0\] _00675_ _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06704_ _02051_ _02186_ _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_07684_ net521 ci_neuron.uut_simple_neuron.titan_id_3\[7\] _03302_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_88_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08686__A1 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04896_ internal_ih.byte4\[4\] _00633_ _00634_ internal_ih.byte0\[4\] _00635_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold442_I internal_ih.byte1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06635_ _01898_ _02274_ _02275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09423_ _04599_ _04650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09354_ _04589_ _04590_ _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06566_ _02166_ _02167_ _02207_ _02208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_75_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08305_ net676 _03821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06497_ _02090_ _02139_ _02140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05517_ _01185_ _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09285_ net85 _04549_ _04552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05448_ _01065_ _01069_ _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08236_ _03748_ _03749_ _03760_ _03747_ _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_132_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08167_ net535 net797 _03702_ _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07118_ _01863_ _02665_ _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05379_ _01049_ _01050_ _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_42_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05424__A1 _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08098_ net548 _00070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07049_ _02555_ _02681_ _02682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_11_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10060_ net197 clknet_leaf_123_sys_clock_i ci_neuron.output_val_internal\[29\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07177__A1 _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07101__A1 _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08601__A1 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10258_ _00551_ clknet_leaf_95_sys_clock_i ci_neuron.stream_o\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05718__A2 _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10189_ _00087_ clknet_leaf_4_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_2\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06420_ _02027_ _02026_ _02064_ _02065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_EDGE_ROW_93_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06351_ _01896_ _01967_ _01996_ _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_84_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06282_ _01878_ _01903_ _01930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05302_ ci_neuron.uut_simple_neuron.x2\[6\] _00861_ _00975_ _00976_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09483__I3 _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09070_ _04378_ net216 _04414_ _00406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05233_ _00863_ _00892_ _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08021_ net607 _00077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold702 ci_neuron.uut_simple_neuron.titan_id_5\[3\] net735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_97_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05164_ _00821_ _00842_ _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold735 _01874_ net768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold724 ci_neuron.input_memory\[1\]\[14\] net804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold713 ci_neuron.uut_simple_neuron.x2\[30\] net746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold746 ci_neuron.uut_simple_neuron.titan_id_5\[31\] net779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout6 net7 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05406__A1 _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold779 ci_neuron.uut_simple_neuron.titan_id_5\[25\] net823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_05095_ _00772_ _00776_ _00777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09972_ _00487_ clknet_leaf_67_sys_clock_i ci_neuron.input_memory\[1\]\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold757 _03544_ net790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold768 ci_neuron.uut_simple_neuron.titan_id_0\[30\] net801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__05618__I _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08923_ _04290_ _04306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08854_ net476 net505 _04264_ _04267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07805_ net602 _00115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05997_ _01611_ _01625_ _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08785_ _04010_ _04211_ _04227_ _00308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04917__B1 _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07736_ ci_neuron.uut_simple_neuron.titan_id_4\[16\] net580 _03345_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04948_ _00666_ _00033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07331__A1 _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07667_ ci_neuron.uut_simple_neuron.titan_id_4\[5\] net629 _03288_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04879_ internal_ih.byte4\[7\] internal_ih.byte3\[7\] _00601_ _00623_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_36_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06618_ _02256_ _02257_ _02258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07598_ _02178_ _03219_ _03222_ _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_94_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09406_ _03742_ net57 _00795_ _01900_ _04622_ _04623_ _04636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_06549_ _02184_ _02190_ _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09337_ _04581_ _00506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09268_ _04138_ _04140_ _04540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07634__A2 _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08219_ _03746_ _00195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09199_ _03742_ _04500_ _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09387__A2 _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10112_ _00236_ clknet_leaf_44_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_4\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_112_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold40 net764 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_54_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10043_ net128 clknet_leaf_113_sys_clock_i ci_neuron.output_val_internal\[12\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold51 ci_neuron.input_memory\[1\]\[11\] net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold62 net809 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold73 _03579_ net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07570__A1 _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold84 internal_ih.spi_tx_byte_o\[2\] net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold95 _00528_ net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07322__A1 _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05920_ _01472_ _01532_ _01579_ _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05851_ _01450_ _01490_ _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer16 _02286_ net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer27 _02938_ net447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08570_ _04052_ _02445_ _04053_ _04054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07521_ _03133_ _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05782_ _01396_ _01399_ _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07452_ _03016_ _03020_ _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08484__I _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07864__A2 ci_neuron.uut_simple_neuron.titan_id_5\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07383_ _03010_ _02859_ _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06403_ _01964_ _02001_ _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_9_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06334_ _01980_ _00169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09122_ _04457_ _00415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08813__A1 _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06265_ _01886_ _01913_ _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09053_ _04383_ net98 ci_neuron.stream_o\[18\] _04384_ _04398_ _04399_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_32_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06196_ _01822_ _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_103_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05216_ ci_neuron.uut_simple_neuron.x2\[0\] _00838_ _00892_ _00893_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_13_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08004_ _03565_ _03567_ _03568_ _03569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold510 ci_neuron.uut_simple_neuron.titan_id_0\[1\] net665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold543 _03369_ net576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05147_ _00824_ _00826_ _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold554 _03648_ net587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold521 net812 net554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold532 _03463_ net565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold565 ci_neuron.uut_simple_neuron.titan_id_3\[9\] net598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold587 ci_neuron.uut_simple_neuron.x0\[13\] net620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold576 _03430_ net609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold598 _03289_ net631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05078_ _00760_ _00757_ _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09955_ _00470_ clknet_leaf_10_sys_clock_i ci_neuron.uut_simple_neuron.x0\[26\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08906_ internal_ih.byte3\[6\] net466 _04296_ _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09886_ _00047_ net19 ci_neuron.value_i\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09392__I2 _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08837_ _04256_ _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_127_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08768_ _00768_ _04214_ _04217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07719_ net457 _00099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08699_ net147 _04136_ _04157_ internal_ih.spi_rx_byte_i\[5\] _04162_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07855__A2 ci_neuron.uut_simple_neuron.titan_id_5\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_138_sys_clock_i clknet_4_2_0_sys_clock_i clknet_leaf_138_sys_clock_i
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_125_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07607__A2 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05094__A2 _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08569__I _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10026_ net92 clknet_leaf_8_sys_clock_i ci_neuron.uut_simple_neuron.titan_id_1\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06346__A2 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07543__A1 ci_neuron.uut_simple_neuron.x3\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09296__A1 _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_3_0_sys_clock_i_I clknet_0_sys_clock_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09048__A1 net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06050_ _00936_ _01706_ _01668_ _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_78_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05001_ _00685_ _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06952_ _02583_ _02586_ _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_94_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09740_ _00319_ clknet_leaf_29_sys_clock_i ci_neuron.uut_simple_neuron.x2\[21\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
.ends

