* NGSPICE file created from ram.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VNW VPW VSS
.ends

.subckt ram address_i[0] address_i[1] address_i[2] address_i[3] address_i[4] clk_i
+ data_i[0] data_i[10] data_i[11] data_i[12] data_i[13] data_i[14] data_i[15] data_i[16]
+ data_i[17] data_i[18] data_i[19] data_i[1] data_i[20] data_i[21] data_i[22] data_i[23]
+ data_i[24] data_i[25] data_i[26] data_i[27] data_i[28] data_i[29] data_i[2] data_i[30]
+ data_i[31] data_i[3] data_i[4] data_i[5] data_i[6] data_i[7] data_i[8] data_i[9]
+ data_o[0] data_o[10] data_o[11] data_o[12] data_o[13] data_o[14] data_o[15] data_o[16]
+ data_o[17] data_o[18] data_o[19] data_o[1] data_o[20] data_o[21] data_o[22] data_o[23]
+ data_o[24] data_o[25] data_o[26] data_o[27] data_o[28] data_o[29] data_o[2] data_o[30]
+ data_o[31] data_o[3] data_o[4] data_o[5] data_o[6] data_o[7] data_o[8] data_o[9]
+ vdd vss we_i
XFILLER_0_118_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5417__B1 _2025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6626__S _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5968__A1 _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7963_ _0263_ clknet_leaf_40_clk_i memory\[20\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4146__S _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6914_ _3434_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7894_ _0194_ clknet_leaf_29_clk_i memory\[18\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_25_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6845_ memory\[14\]\[0\] _1164_ _3397_ _3398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_135_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6776_ _3360_ _3361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_17_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3988_ net25 _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6393__A1 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8515_ _0815_ clknet_leaf_118_clk_i memory\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5727_ _1957_ memory\[26\]\[9\] _2335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_115_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8446_ _0746_ clknet_leaf_198_clk_i memory\[13\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5658_ _1988_ memory\[0\]\[7\] _2268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6940__I0 _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7192__S _3578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5589_ _1856_ _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4609_ memory\[21\]\[28\] _1229_ _1509_ _1518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8377_ _0677_ clknet_leaf_0_clk_i memory\[14\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7328_ _1104_ memory\[4\]\[3\] _3650_ _3654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7259_ _3617_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_5_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5959__A1 _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4482__I1 _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3895__S _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5615__S _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6931__I0 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6687__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__I _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3869__I net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4960_ _1089_ memory\[26\]\[30\] _1673_ _1707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7277__S _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3911_ net28 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_59_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ _1670_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6375__A1 _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6630_ _1987_ memory\[11\]\[28\] _3218_ _1907_ _3219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_104_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6561_ _2796_ net57 _3152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8300_ _0600_ clknet_leaf_58_clk_i net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_133_clk_i_I clknet_4_9_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5512_ memory\[12\]\[4\] memory\[13\]\[4\] _1978_ _2125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6492_ _3081_ _2760_ _3083_ _2716_ _3084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_70_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8231_ _0531_ clknet_leaf_114_clk_i memory\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5443_ memory\[24\]\[3\] _1859_ _2057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5374_ _1872_ _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8162_ _0462_ clknet_leaf_165_clk_i memory\[27\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7113_ _3539_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4325_ _1364_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5324__I _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8093_ _0393_ clknet_leaf_8_clk_i memory\[24\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4256_ _1078_ memory\[29\]\[25\] _1322_ _1328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7044_ _3502_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4161__I0 _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6356__S _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4187_ _1288_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_58_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6155__I _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7946_ _0246_ clknet_leaf_131_clk_i memory\[20\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7877_ _0177_ clknet_leaf_143_clk_i memory\[18\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6091__S _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5927__C _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5169__A2 _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6828_ _3388_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6759_ _3342_ _3344_ _1890_ _3345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6118__A1 _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8429_ _0729_ clknet_leaf_64_clk_i memory\[13\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6913__I0 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6669__A2 _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4152__I0 _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6065__I _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7641__I1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6357__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4313__I _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7560__S _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5144__I _1782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4110_ _1238_ _1062_ _1166_ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5090_ _1776_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4143__I0 _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4041_ _1170_ _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5992_ _2310_ memory\[11\]\[14\] _2594_ _2174_ _2595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7632__I1 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7800_ _0100_ clknet_leaf_220_clk_i memory\[15\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7731_ _0031_ clknet_leaf_31_clk_i memory\[19\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4943_ _1698_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5747__C _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7662_ _3830_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4874_ _1070_ memory\[25\]\[21\] _1660_ _1662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7396__I0 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6613_ _1932_ _3201_ _1856_ _3202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7593_ _3757_ _1522_ _3794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_43_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6544_ _3132_ _2872_ _3134_ _2826_ _3135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__5763__B _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6475_ _2933_ _3064_ _3066_ _3067_ _3068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_8214_ _0514_ clknet_leaf_14_clk_i memory\[28\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5426_ _2038_ _2040_ _1939_ _2041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6578__C _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7470__S _3722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8145_ _0445_ clknet_leaf_43_clk_i memory\[26\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5357_ memory\[16\]\[1\] memory\[17\]\[1\] _1911_ _1973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8076_ _0376_ clknet_leaf_55_clk_i memory\[24\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4308_ _1355_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5288_ _1863_ _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6086__S _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input36_I data_i[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4239_ _1275_ memory\[29\]\[17\] _1311_ _1319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7027_ memory\[13\]\[22\] _1217_ _3491_ _3494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6814__S _3372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6587__A1 _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7929_ _0229_ clknet_leaf_208_clk_i memory\[1\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4334__S _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7645__S _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_137_Right_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5165__S _1782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6511__A1 _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4373__I0 _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7380__S _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4509__S _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4676__I1 _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6578__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7378__I0 _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4590_ memory\[21\]\[19\] _1210_ _1498_ _1508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6679__B _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6260_ memory\[30\]\[20\] memory\[31\]\[20\] _2532_ _2857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_110_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6191_ memory\[4\]\[18\] _2468_ _2790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5211_ _1840_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5142_ _1137_ memory\[2\]\[19\] _1794_ _1804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7302__I0 _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _1767_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4419__S _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4024_ _1180_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7605__I1 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6569__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5758__B _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ _2288_ _2577_ _2200_ _2578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4926_ _1689_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7714_ _0014_ clknet_leaf_137_clk_i memory\[19\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5477__C _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8694_ _0994_ clknet_leaf_191_clk_i memory\[5\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4857_ _1267_ memory\[25\]\[13\] _1649_ _1653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7645_ memory\[6\]\[24\] net22 _3817_ _3822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7576_ _3785_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4788_ _1616_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6527_ _2000_ memory\[29\]\[26\] _3117_ _2855_ _3118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_95_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6458_ memory\[12\]\[24\] memory\[13\]\[24\] _2919_ _3051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5409_ memory\[23\]\[2\] _1896_ _2023_ _1899_ _2024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6389_ _2981_ memory\[7\]\[22\] _2982_ _2983_ _2984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__3858__A2 _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8128_ _0428_ clknet_leaf_133_clk_i memory\[25\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8059_ _0359_ clknet_leaf_11_clk_i memory\[23\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3967__I _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6343__I _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6732__A1 _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4346__I0 _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5850__C _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4649__I1 _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4239__S _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5471__A1 _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5774__A2 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5760_ _2318_ memory\[0\]\[9\] _2368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6253__I _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4711_ _1260_ memory\[23\]\[10\] _1573_ _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5691_ memory\[16\]\[8\] memory\[17\]\[8\] _2164_ _2300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7285__S _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4642_ _1536_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7430_ _3707_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4702__S _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5526__A2 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4573_ _1499_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7361_ _1137_ memory\[4\]\[19\] _3661_ _3671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7292_ _3634_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6312_ memory\[22\]\[21\] _2908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6243_ _2515_ memory\[7\]\[19\] _2840_ _2517_ _2841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_12_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6174_ _1879_ _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4149__S _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5125_ _1795_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5056_ _1260_ memory\[28\]\[10\] _1758_ _1759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4007_ _1059_ _1060_ _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5462__A1 _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5765__A2 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8746_ _1046_ clknet_leaf_85_clk_i memory\[7\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5958_ _1863_ _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4812__I1 _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4909_ _1680_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5889_ memory\[16\]\[12\] memory\[17\]\[12\] _2164_ _2494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8677_ _0977_ clknet_leaf_119_clk_i memory\[5\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5935__C _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7628_ memory\[6\]\[16\] net13 _3806_ _3813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_97_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_181_clk_i_I clknet_4_9_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6714__A1 _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7559_ _3776_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7514__I0 _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5951__B _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4328__I0 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6338__I _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5242__I _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3898__S _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__I _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5845__C _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5692__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5444__A1 _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6930_ _3442_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6861_ memory\[14\]\[8\] _1187_ _3397_ _3406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5812_ memory\[2\]\[10\] memory\[3\]\[10\] _2270_ _2419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6792_ _3369_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8600_ _0900_ clknet_leaf_210_clk_i memory\[4\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5743_ _2160_ memory\[19\]\[9\] _2350_ _2075_ _2351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8531_ _0831_ clknet_leaf_83_clk_i memory\[8\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8462_ _0762_ clknet_leaf_60_clk_i memory\[31\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5674_ _1862_ memory\[27\]\[8\] _2282_ _1867_ _2283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_7413_ _1121_ memory\[0\]\[11\] _3697_ _3699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8393_ _0693_ clknet_leaf_125_clk_i memory\[16\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_79_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4625_ _1527_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7344_ _3662_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4556_ _1490_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7275_ _1118_ memory\[3\]\[10\] _3625_ _3626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_92_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4487_ _1453_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6586__C _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6226_ memory\[12\]\[19\] memory\[13\]\[19\] _2453_ _2824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6158__I _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6157_ _2754_ _2755_ _2666_ _2756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_128_clk_i_I clknet_4_14_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5108_ _1786_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6088_ _2686_ _2688_ _2414_ _2689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5435__A1 _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4607__S _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5039_ _1244_ memory\[28\]\[2\] _1747_ _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4410__A2 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8729_ _1029_ clknet_leaf_1_clk_i memory\[6\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_134_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6163__A2 _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4141__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5237__I net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7653__S _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5681__B _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput42 net42 data_o[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5173__S _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6269__S _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput64 net64 data_o[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput53 net53 data_o[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4721__I0 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5674__A1 _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4517__S _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5029__I1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5348__S _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5575__C _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4252__S _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4410_ _1057_ net4 _1063_ _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__5591__B _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5390_ _1371_ _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_23_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4341_ _1373_ _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5083__S _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4960__I0 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3890__I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7060_ memory\[31\]\[5\] _1181_ _3506_ _3512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_74_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4272_ _1237_ memory\[17\]\[0\] _1336_ _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5665__A1 _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6011_ _2432_ memory\[26\]\[15\] _2613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_94_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6907__S _3396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4427__S _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7962_ _0262_ clknet_leaf_39_clk_i memory\[20\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6090__A1 _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6913_ _1093_ memory\[16\]\[0\] _3433_ _3434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_12_0_clk_i clknet_0_clk_i clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7893_ _0193_ clknet_leaf_27_clk_i memory\[18\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6844_ _3396_ _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6775_ _1298_ _3359_ _3360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3987_ _1153_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6393__A2 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5726_ memory\[24\]\[9\] _2333_ _2334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8514_ _0814_ clknet_leaf_146_clk_i memory\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8445_ _0745_ clknet_leaf_216_clk_i memory\[13\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_54_clk_i_I clknet_4_5_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6145__A2 _2732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5657_ _1903_ _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5588_ memory\[30\]\[6\] memory\[31\]\[6\] _2066_ _2199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4608_ _1517_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8376_ _0676_ clknet_leaf_0_clk_i memory\[14\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4539_ _1480_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7327_ _3653_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3903__A1 _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7258_ _1102_ memory\[3\]\[2\] _3614_ _3617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6209_ _2529_ memory\[29\]\[19\] _2806_ _2389_ _2807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_7189_ _3580_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_5_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6552__S _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_172_clk_i clknet_4_8_0_clk_i clknet_leaf_172_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_106_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_187_clk_i clknet_4_3_0_clk_i clknet_leaf_187_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_114_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4942__I0 _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Left_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_39_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_110_clk_i clknet_4_15_0_clk_i clknet_leaf_110_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5647__A1 _2240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_125_clk_i clknet_4_14_0_clk_i clknet_leaf_125_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7558__S _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_129_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4890_ _1086_ memory\[25\]\[29\] _1660_ _1670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3910_ _1101_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6560_ _3135_ _3140_ _3145_ _3150_ _2894_ _3151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_82_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5511_ memory\[14\]\[4\] _2124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6127__A2 _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7293__S _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6491_ memory\[23\]\[25\] _2713_ _3082_ _2671_ _3083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_54_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8230_ _0530_ clknet_leaf_116_clk_i memory\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_57_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5442_ _1855_ _2032_ _2055_ _2056_ _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_30_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4933__I0 _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5373_ _1988_ memory\[0\]\[1\] _1989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_10_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8161_ _0461_ clknet_leaf_174_clk_i memory\[27\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8092_ _0392_ clknet_leaf_7_clk_i memory\[24\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7112_ memory\[31\]\[30\] _1233_ _3505_ _3539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4324_ _1078_ memory\[17\]\[25\] _1358_ _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7043_ memory\[13\]\[30\] _1233_ _3468_ _3502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5541__S _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4255_ _1327_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4186_ _1082_ memory\[15\]\[27\] _1280_ _1288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_2_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6063__A1 _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6989__I1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5810__A1 _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7468__S _3722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7945_ _0245_ clknet_leaf_129_clk_i memory\[20\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7876_ _0176_ clknet_leaf_142_clk_i memory\[18\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6827_ _1148_ memory\[9\]\[24\] _3383_ _3388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_108_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6104__C _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6758_ _1909_ _3343_ _1994_ _3344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5709_ _1869_ _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6689_ memory\[24\]\[30\] _1858_ _3276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7166__I1 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8428_ _0728_ clknet_leaf_61_clk_i memory\[13\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5177__I0 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4620__S _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5877__A1 _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8359_ _0659_ clknet_leaf_150_clk_i memory\[14\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5629__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6547__S _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_42_clk_i clknet_4_4_0_clk_i clknet_leaf_42_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5250__I _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7378__S _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_57_clk_i clknet_4_7_0_clk_i clknet_leaf_57_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5801__B2 _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7157__I1 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4530__S _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__A1 _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6030__B _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4040_ net7 _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6293__A1 _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6045__A1 _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5991_ _2362_ memory\[10\]\[14\] _2594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7730_ _0030_ clknet_leaf_74_clk_i memory\[19\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4942_ _1070_ memory\[26\]\[21\] _1696_ _1698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7661_ _1093_ memory\[7\]\[0\] _1087_ _3830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_35_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4873_ _1661_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6612_ memory\[30\]\[28\] memory\[31\]\[28\] _1923_ _3201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5556__B1 _2159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7592_ _3793_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_65_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6543_ memory\[15\]\[26\] _2823_ _3133_ _2773_ _3134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_40_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4440__S _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__I0 _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6474_ _2938_ _2939_ memory\[5\]\[24\] _3067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5859__A1 _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5425_ _1934_ _2039_ _1937_ _2040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8213_ _0513_ clknet_leaf_23_clk_i memory\[28\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4906__I0 _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5335__I _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8144_ _0444_ clknet_leaf_48_clk_i memory\[26\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5356_ _1904_ memory\[19\]\[1\] _1971_ _1907_ _1972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4307_ _1275_ memory\[17\]\[17\] _1347_ _1355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8075_ _0375_ clknet_leaf_45_clk_i memory\[24\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5287_ _1903_ _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_10_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4238_ _1318_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_74_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7026_ _3493_ _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input29_I data_i[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4169_ _1056_ memory\[15\]\[19\] _1261_ _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7198__S _3578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5938__C _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4615__S _1486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6831__I0 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7928_ _0228_ clknet_leaf_193_clk_i memory\[1\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7859_ _0159_ clknet_leaf_32_clk_i memory\[17\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6339__A2 _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_83_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7139__I1 _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4350__S _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7661__S _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5245__I _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_92_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5181__S _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_176_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4260__S _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5583__C _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7550__I1 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5210_ _1137_ memory\[30\]\[19\] _1830_ _1840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6502__A2 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7571__S _3781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6190_ _2786_ _2788_ _2421_ _2789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5141_ _1803_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5091__S _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5072_ _1277_ memory\[28\]\[18\] _1758_ _1767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4023_ memory\[12\]\[4\] _1179_ _1171_ _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6018__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6915__S _3433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5974_ memory\[30\]\[14\] memory\[31\]\[14\] _2532_ _2577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7713_ _0013_ clknet_leaf_178_clk_i memory\[19\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4925_ _1267_ memory\[26\]\[13\] _1685_ _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8693_ _0993_ clknet_leaf_187_clk_i memory\[5\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4856_ _1652_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7644_ _3821_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7575_ memory\[5\]\[23\] net21 _3781_ _3785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4787_ memory\[24\]\[12\] _1196_ _1613_ _1616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6526_ _2001_ memory\[28\]\[26\] _3117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_43_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7481__S _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7541__I1 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6457_ memory\[14\]\[24\] _3050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_100_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5408_ memory\[20\]\[2\] memory\[21\]\[2\] _1897_ _2023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6388_ _1866_ _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8127_ _0427_ clknet_leaf_183_clk_i memory\[25\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5339_ _1855_ _1919_ _1953_ _1955_ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6257__A1 _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8058_ _0358_ clknet_leaf_11_clk_i memory\[23\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7009_ _3484_ _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6009__A1 _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6825__S _3383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6804__I0 _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6496__A1 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6248__A1 _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7296__I0 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5859__B _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5578__C _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6420__A1 _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7566__S _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4282__I0 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5690_ _2160_ memory\[19\]\[8\] _2298_ _2075_ _2299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4710_ _1561_ _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_57_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4641_ memory\[22\]\[10\] _1191_ _1535_ _1536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6723__A2 _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4572_ memory\[21\]\[10\] _1191_ _1498_ _1499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7360_ _3670_ _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7291_ _1135_ memory\[3\]\[18\] _3625_ _3634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6311_ _2904_ _2906_ _2757_ _2907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_122_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6242_ _2562_ memory\[6\]\[19\] _2840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6487__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7287__I0 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6239__A1 _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6173_ memory\[12\]\[18\] memory\[13\]\[18\] _2453_ _2772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5124_ _1260_ memory\[2\]\[10\] _1794_ _1795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5055_ _1746_ _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4006_ _1057_ _1166_ _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_95_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ memory\[4\]\[13\] _2468_ _2561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8745_ _1045_ clknet_leaf_104_clk_i memory\[7\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7476__S _3722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8676_ _0976_ clknet_leaf_118_clk_i memory\[5\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4908_ _1250_ memory\[26\]\[5\] _1674_ _1680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7211__I0 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7627_ _3812_ _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5888_ _2160_ memory\[19\]\[12\] _2492_ _2075_ _2493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_63_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_124_clk_i_I clknet_4_14_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4839_ _1643_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4576__I1 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7558_ memory\[5\]\[15\] net12 _3770_ _3776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7489_ _1129_ memory\[10\]\[15\] _3733_ _3739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6509_ _2733_ memory\[1\]\[25\] _3100_ _2975_ _3101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_132_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5523__I _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_49_clk_i_I clknet_4_5_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4500__I1 _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6650__A1 _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_11_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4264__I0 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7450__I0 _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4964__A1 _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7386__S _3649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7202__I0 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7185__I _3577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4567__I1 _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_20_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_117_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6469__A1 _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6641__A1 _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6860_ _3405_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6791_ _1112_ memory\[9\]\[7\] _3361_ _3369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5811_ _1882_ _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8530_ _0830_ clknet_leaf_95_clk_i memory\[8\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4713__S _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5742_ _2208_ memory\[18\]\[9\] _2350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_91_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7296__S _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8461_ _0761_ clknet_leaf_60_clk_i memory\[31\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5673_ _1957_ memory\[26\]\[8\] _2282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7412_ _3698_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8392_ _0692_ clknet_leaf_111_clk_i memory\[16\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4624_ memory\[22\]\[2\] _1175_ _1524_ _1527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7343_ _1118_ memory\[4\]\[10\] _3661_ _3662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4555_ memory\[21\]\[2\] _1175_ _1487_ _1490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7274_ _3613_ _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4486_ memory\[20\]\[2\] _1175_ _1450_ _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6225_ _1895_ _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6156_ memory\[30\]\[18\] memory\[31\]\[18\] _2532_ _2755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5107_ _1244_ memory\[2\]\[2\] _1783_ _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6087_ _2313_ _2687_ _2643_ _2688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_50_clk_i_I clknet_4_5_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7680__I0 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5499__B _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6632__A1 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input11_I data_i[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5038_ _1749_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6174__I _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4246__I0 _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7432__I0 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6989_ memory\[13\]\[4\] _1179_ _3469_ _3474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8728_ _1028_ clknet_leaf_1_clk_i memory\[6\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5946__C _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4797__I1 _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4410__A3 _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8659_ _0959_ clknet_leaf_77_clk_i memory\[10\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput43 net43 data_o[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_102_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput65 net65 data_o[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5253__I _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput54 net54 data_o[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__7671__I0 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7423__I0 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4237__I0 _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5428__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4340_ net38 _1372_ _1373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_10_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4271_ _1335_ _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6010_ memory\[24\]\[15\] _2333_ _2612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input3_I address_i[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4708__S _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7961_ _0261_ clknet_leaf_40_clk_i memory\[20\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6923__S _3433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6912_ _3432_ _3433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7892_ _0192_ clknet_leaf_28_clk_i memory\[18\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6843_ _1167_ _1522_ _3396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_76_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6774_ _1057_ _3358_ _3359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3986_ memory\[19\]\[26\] _1152_ _1140_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5725_ _1858_ _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_73_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8513_ _0813_ clknet_leaf_147_clk_i memory\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5656_ _2263_ _2265_ _1939_ _2266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8444_ _0744_ clknet_leaf_218_clk_i memory\[13\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4607_ memory\[21\]\[27\] _1227_ _1509_ _1517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5587_ _2063_ memory\[29\]\[6\] _2197_ _1880_ _2198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4400__I0 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5353__B2 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8375_ _0675_ clknet_leaf_220_clk_i memory\[14\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7326_ _1102_ memory\[4\]\[2\] _3650_ _3653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4538_ memory\[20\]\[27\] _1227_ _1472_ _1480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6169__I _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7257_ _3616_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4469_ _1082_ memory\[1\]\[27\] _1435_ _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6208_ _2574_ memory\[28\]\[19\] _2806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7188_ _1100_ memory\[8\]\[1\] _3578_ _3580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6139_ _2735_ _2738_ _2421_ _2739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_5_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4467__I0 _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6833__S _3383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6369__B1 _2957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5692__B _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3991__I net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5344__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4528__S _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__A2 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_103_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5583__A1 _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4062__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5510_ _2107_ _2113_ _2117_ _2122_ _1918_ _2123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_55_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6490_ memory\[20\]\[25\] memory\[21\]\[25\] _2812_ _3082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6698__B _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5441_ _1954_ net61 _2056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5886__A2 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_112_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5372_ _1869_ _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8160_ _0460_ clknet_leaf_135_clk_i memory\[26\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4323_ _1363_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8091_ _0391_ clknet_leaf_7_clk_i memory\[24\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7111_ _3538_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7042_ _3501_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4254_ _1076_ memory\[29\]\[24\] _1322_ _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4438__S _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4185_ _1287_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7944_ _0244_ clknet_leaf_153_clk_i memory\[20\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5269__S _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7875_ _0175_ clknet_leaf_138_clk_i memory\[18\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6826_ _3387_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5574__A1 _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6757_ memory\[8\]\[31\] memory\[9\]\[31\] _1992_ _3343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5708_ _2312_ _2316_ _1939_ _2317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_70_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3969_ _1141_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6688_ _2846_ _3254_ _3274_ _3275_ _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_104_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8427_ _0727_ clknet_leaf_77_clk_i memory\[13\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5639_ memory\[23\]\[7\] _2247_ _2248_ _2205_ _2249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_131_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8358_ _0658_ clknet_leaf_157_clk_i memory\[14\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7309_ _3643_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8289_ _0589_ clknet_leaf_140_clk_i net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5629__A2 _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4348__S _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output42_I net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7659__S _3794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5801__A2 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5179__S _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7394__S _3686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_172_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6311__B _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__A2 _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6738__S _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4258__S _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7569__S _3781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_97_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5990_ _2590_ _2406_ _2592_ _2360_ _2593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__4851__I0 _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4941_ _1697_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5089__S _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4872_ _1068_ memory\[25\]\[20\] _1660_ _1661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6272__I _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7660_ _3829_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5556__A1 _2150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6611_ _2000_ memory\[29\]\[28\] _3199_ _2855_ _3200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_90_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7591_ memory\[5\]\[31\] net30 _3758_ _3793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4721__S _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6542_ memory\[12\]\[26\] memory\[13\]\[26\] _2919_ _3133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6221__B _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6473_ _2981_ memory\[7\]\[24\] _3065_ _2983_ _3066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8212_ _0512_ clknet_leaf_34_clk_i memory\[28\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5424_ memory\[8\]\[2\] memory\[9\]\[2\] _1935_ _2039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8143_ _0443_ clknet_leaf_48_clk_i memory\[26\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6520__A3 _3110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5355_ _1905_ memory\[18\]\[1\] _1971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4306_ _1354_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8074_ _0374_ clknet_leaf_130_clk_i memory\[24\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5286_ _1295_ _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_10_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4237_ _1273_ memory\[29\]\[16\] _1311_ _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_171_clk_i clknet_4_8_0_clk_i clknet_leaf_171_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7025_ memory\[13\]\[21\] _1215_ _3491_ _3493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6036__A2 _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7479__S _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4168_ _1278_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5095__I0 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4099_ net27 _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_78_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_186_clk_i clknet_4_3_0_clk_i clknet_leaf_186_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4842__I0 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7927_ _0227_ clknet_leaf_193_clk_i memory\[1\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7858_ _0158_ clknet_leaf_74_clk_i memory\[17\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5300__B _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6809_ _3378_ _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7789_ _0089_ clknet_leaf_63_clk_i memory\[15\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6131__B _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_124_clk_i clknet_4_14_0_clk_i clknet_leaf_124_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_14_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_139_clk_i clknet_4_10_0_clk_i clknet_leaf_139_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_119_clk_i_I clknet_4_14_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7075__I1 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4806__S _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5538__A1 _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5436__I _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6889__I1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5710__A1 _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6695__C _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6468__S _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5140_ _1277_ memory\[2\]\[18\] _1794_ _1803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5071_ _1766_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6266__A2 _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4022_ net32 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7066__I1 _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5077__I0 _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5973_ _2529_ memory\[29\]\[14\] _2575_ _2389_ _2576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_84_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4924_ _1688_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6931__S _3433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7712_ _0012_ clknet_leaf_179_clk_i memory\[7\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8692_ _0992_ clknet_leaf_79_clk_i memory\[5\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4855_ _1265_ memory\[25\]\[12\] _1649_ _1652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5529__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7643_ memory\[6\]\[23\] net21 _3817_ _3821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4786_ _1615_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7574_ _3784_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_41_clk_i clknet_4_4_0_clk_i clknet_leaf_41_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6525_ _2798_ _3112_ _3114_ _3115_ _3116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_16_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ _3034_ _3039_ _3043_ _3048_ _2869_ _3049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_3_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5407_ memory\[22\]\[2\] _2022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6387_ _2562_ memory\[6\]\[22\] _2982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_56_clk_i clknet_4_5_0_clk_i clknet_leaf_56_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_101_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8126_ _0426_ clknet_leaf_17_clk_i memory\[25\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5338_ _1954_ net39 _1955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6177__I _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8057_ _0357_ clknet_leaf_39_clk_i memory\[23\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7008_ memory\[13\]\[13\] _1198_ _3480_ _3484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_126_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_120_clk_i_I clknet_4_14_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5269_ memory\[30\]\[0\] memory\[31\]\[0\] _1885_ _1886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7002__S _3480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5068__I0 _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4626__S _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5768__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6841__S _3360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5457__S _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6193__A1 _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5940__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4160__I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_45_clk_i_I clknet_4_5_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5256__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5192__S _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6288__S _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4536__S _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4640_ _1523_ _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_71_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5231__I0 _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4571_ _1486_ _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_71_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6310_ _2754_ _2905_ _2666_ _2906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7290_ _3633_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6241_ memory\[4\]\[19\] _2468_ _2839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6172_ memory\[14\]\[18\] _2771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5123_ _1782_ _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5054_ _1757_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4446__S _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4005_ _1165_ _1063_ _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__7039__I1 _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6798__I0 _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4245__I _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5956_ _2557_ _2559_ _2421_ _2560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8744_ _1044_ clknet_leaf_109_clk_i memory\[7\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5887_ _2208_ memory\[18\]\[12\] _2492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5785__B _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8675_ _0975_ clknet_leaf_144_clk_i memory\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4907_ _1679_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7626_ memory\[6\]\[15\] net12 _3806_ _3812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4838_ _1248_ memory\[25\]\[4\] _1638_ _1643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6175__B2 _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7557_ _3775_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5076__I _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4769_ _1606_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7488_ _3738_ _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6508_ _2784_ memory\[0\]\[25\] _3100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_132_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6439_ _2848_ memory\[27\]\[24\] _3031_ _2850_ _3032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_132_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8109_ _0409_ clknet_leaf_56_clk_i memory\[25\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_54_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5989__B2 _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4356__S _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6650__A2 _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6789__I0 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7667__S _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_65_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3994__I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6166__A1 _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5187__S _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4091__S _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5213__I0 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5913__A1 _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6961__I0 _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4266__S _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7577__S _3781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5810_ _2267_ memory\[1\]\[10\] _2416_ _2043_ _2417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6790_ _3368_ _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4065__I net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5741_ _2345_ _2294_ _2348_ _2250_ _2349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_18_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8460_ _0760_ clknet_leaf_59_clk_i memory\[31\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5097__S _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5204__I0 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7411_ _1118_ memory\[0\]\[10\] _3697_ _3698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6157__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5672_ memory\[24\]\[8\] _1859_ _2281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8391_ _0691_ clknet_leaf_124_clk_i memory\[16\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6952__I0 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4623_ _1526_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7342_ _3649_ _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4554_ _1489_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7273_ _3624_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6224_ memory\[14\]\[19\] _2822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4485_ _1452_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6155_ _1882_ _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6086_ memory\[8\]\[16\] memory\[9\]\[16\] _2314_ _2687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5106_ _1785_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5037_ _1242_ memory\[28\]\[1\] _1747_ _1749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4176__S _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4494__I1 _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7487__S _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6396__A1 _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4904__S _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6988_ _3473_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8727_ _1027_ clknet_leaf_192_clk_i memory\[6\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5939_ memory\[16\]\[13\] memory\[17\]\[13\] _2164_ _2543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_101_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6404__B _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8658_ _0958_ clknet_leaf_65_clk_i memory\[10\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7196__I0 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6123__C _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_218_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8589_ _0889_ clknet_leaf_93_clk_i memory\[4\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7609_ memory\[6\]\[7\] net35 _3795_ _3803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput44 net44 data_o[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput66 net66 data_o[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput55 net55 data_o[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_101_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4182__I0 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4814__S _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6387__A1 _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5709__I _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_119_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6934__I0 _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ _1095_ _1298_ _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_94_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6275__I _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5822__B1 _2422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7960_ _0260_ clknet_leaf_40_clk_i memory\[20\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_167_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7891_ _0191_ clknet_leaf_31_clk_i memory\[18\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6911_ _1095_ _1598_ _3432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6842_ _3395_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7100__S _3528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4523__I _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6773_ net4 _1094_ _3358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_18_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3985_ net24 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_116_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5724_ _1856_ _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8512_ _0812_ clknet_leaf_174_clk_i memory\[11\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6925__I0 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5655_ _1934_ _2264_ _2177_ _2265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8443_ _0743_ clknet_leaf_217_clk_i memory\[13\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4606_ _1516_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8374_ _0674_ clknet_leaf_5_clk_i memory\[14\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5586_ _2108_ memory\[28\]\[6\] _2197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7325_ _3652_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6550__A1 _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5353__A2 _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4537_ _1479_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7256_ _1100_ memory\[3\]\[1\] _3614_ _3616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4468_ _1442_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4164__I0 _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6207_ _2798_ _2800_ _2802_ _2804_ _2805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_68_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7187_ _3579_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6138_ _2418_ _2737_ _2602_ _2738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4399_ _1405_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6185__I _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ memory\[20\]\[16\] memory\[21\]\[16\] _2346_ _2670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_6_0_clk_i clknet_0_clk_i clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6605__A2 _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7653__I1 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4634__S _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6369__A1 _2948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7010__S _3480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4433__I _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5344__A2 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7680__S _3837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4155__I0 _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4544__S _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4343__I _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4630__I1 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_132_Right_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ _2036_ _2041_ _2047_ _2054_ _1952_ _2055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_42_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_93_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5371_ _1903_ _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4394__I0 _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7332__I0 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4322_ _1076_ memory\[17\]\[24\] _1358_ _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8090_ _0390_ clknet_leaf_8_clk_i memory\[24\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7110_ memory\[31\]\[29\] _1231_ _3528_ _3538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4146__I0 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4719__S _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4253_ _1326_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7041_ memory\[13\]\[29\] _1231_ _3491_ _3501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4184_ _1080_ memory\[15\]\[26\] _1280_ _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6934__S _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6599__A1 _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7943_ _0243_ clknet_leaf_155_clk_i memory\[20\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5271__A1 _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7874_ _0174_ clknet_leaf_138_clk_i memory\[18\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6825_ _1146_ memory\[9\]\[23\] _3383_ _3387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_135_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3968_ memory\[19\]\[20\] _1139_ _1140_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6771__A1 _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6756_ _1987_ memory\[11\]\[31\] _3341_ _1907_ _3342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5707_ _2313_ _2315_ _2177_ _2316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_72_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6687_ _1854_ net60 _3275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3899_ _1092_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_131_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6401__C _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5326__A2 _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5638_ memory\[20\]\[7\] memory\[21\]\[7\] _1897_ _2248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8426_ _0726_ clknet_leaf_178_clk_i memory\[13\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6523__A1 _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5569_ _1987_ memory\[1\]\[5\] _2180_ _2043_ _2181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_13_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8357_ _0657_ clknet_leaf_157_clk_i memory\[14\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7308_ _1152_ memory\[3\]\[26\] _3636_ _3643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8288_ _0588_ clknet_leaf_180_clk_i memory\[30\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_129_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7239_ _3606_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_129_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7626__I1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5259__I _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4163__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_115_clk_i_I clknet_4_15_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_1_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6514__A1 _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7314__I0 _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4828__A1 _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6818__I _3360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4338__I _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4940_ _1068_ memory\[26\]\[20\] _1696_ _1697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4274__S _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4871_ _1637_ _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6610_ _2001_ memory\[28\]\[28\] _3199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7585__S _3781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7590_ _3792_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4603__I1 _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6541_ memory\[14\]\[26\] _3132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6753__B2 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6472_ _1864_ memory\[6\]\[24\] _3065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4367__I0 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6929__S _3433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8211_ _0511_ clknet_leaf_34_clk_i memory\[28\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5423_ _1929_ memory\[11\]\[2\] _2037_ _1932_ _2038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_11_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5833__S _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8142_ _0442_ clknet_leaf_47_clk_i memory\[26\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5354_ _1967_ _1894_ _1969_ _1901_ _1970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4305_ _1273_ memory\[17\]\[16\] _1347_ _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5285_ _1892_ _1894_ _1900_ _1901_ _1902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_8073_ _0373_ clknet_leaf_177_clk_i memory\[24\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4236_ _1317_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7024_ _3492_ _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4167_ _1277_ memory\[15\]\[18\] _1261_ _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5492__A1 _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4098_ _1230_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4184__S _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7926_ _0226_ clknet_leaf_194_clk_i memory\[1\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7857_ _0157_ clknet_leaf_71_clk_i memory\[17\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6808_ _1129_ memory\[9\]\[15\] _3372_ _3378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7495__S _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4912__S _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7788_ _0088_ clknet_leaf_61_clk_i memory\[15\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5547__A2 _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5807__I _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _1932_ _3324_ _1856_ _3325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6412__B _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4358__I0 _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8409_ _0709_ clknet_leaf_20_clk_i memory\[16\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6839__S _3360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_131_Left_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5483__A1 _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6574__S _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_41_clk_i_I clknet_4_4_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3997__I net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4094__S _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4822__S _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6735__A1 _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5452__I _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5070_ _1275_ memory\[28\]\[17\] _1758_ _1766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4068__I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5474__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4021_ _1178_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5972_ _2574_ memory\[28\]\[14\] _2575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6283__I _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4923_ _1265_ memory\[26\]\[12\] _1685_ _1688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__I1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7711_ _0011_ clknet_leaf_179_clk_i memory\[7\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8691_ _0991_ clknet_leaf_78_clk_i memory\[5\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4732__S _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4854_ _1651_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5529__A2 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6726__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7642_ _3820_ _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4785_ memory\[24\]\[11\] _1194_ _1613_ _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7573_ memory\[5\]\[22\] net20 _3781_ _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6524_ _2803_ _1990_ memory\[25\]\[26\] _3115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_43_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6455_ _3045_ _3047_ _2768_ _3048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_42_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5790__C _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5406_ _2018_ _2020_ _1890_ _2021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6386_ _1861_ _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_100_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8125_ _0425_ clknet_leaf_4_clk_i memory\[25\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5337_ _1854_ _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5362__I _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8056_ _0356_ clknet_leaf_40_clk_i memory\[23\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5268_ _1884_ _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7007_ _3483_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_126_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input34_I data_i[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4219_ _1308_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5199_ _1834_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6009__A3 _2610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5768__A2 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6414__B1 _3002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7909_ _0209_ clknet_leaf_119_clk_i memory\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_137_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5473__S _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6248__A3 _2844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6036__C _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4806__I1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5875__C _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4570_ _1497_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_170_clk_i clknet_4_8_0_clk_i clknet_leaf_170_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5891__B _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7508__I0 _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6240_ _2835_ _2837_ _2421_ _2838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_94_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6171_ _2751_ _2758_ _2763_ _2769_ _2403_ _2770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5695__A1 _2285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4742__I0 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_185_clk_i clknet_4_3_0_clk_i clknet_leaf_185_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ _1793_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5447__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5910__I _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5053_ _1258_ memory\[28\]\[9\] _1747_ _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4727__S _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4004_ net4 _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__6942__S _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_123_clk_i clknet_4_14_0_clk_i clknet_leaf_123_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5955_ _2418_ _2558_ _2136_ _2559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8743_ _1043_ clknet_leaf_107_clk_i memory\[7\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5558__S _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5886_ _2488_ _2294_ _2490_ _2250_ _2491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_118_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8674_ _0974_ clknet_leaf_144_clk_i memory\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4906_ _1248_ memory\[26\]\[4\] _1674_ _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7625_ _3811_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_106_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4837_ _1642_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6175__A2 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_138_clk_i clknet_4_9_0_clk_i clknet_leaf_138_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7556_ memory\[5\]\[14\] net11 _3770_ _3775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_9_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4768_ memory\[24\]\[3\] _1177_ _1602_ _1606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7487_ _1127_ memory\[10\]\[14\] _3733_ _3738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6507_ _3096_ _3098_ _2880_ _3099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_16_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4699_ _1567_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6438_ _2898_ memory\[26\]\[24\] _3031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_132_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8108_ _0408_ clknet_leaf_46_clk_i memory\[25\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6369_ _2948_ _2953_ _2957_ _2963_ _2869_ _2964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5438__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_214_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5989__A2 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8039_ _0339_ clknet_leaf_154_clk_i memory\[23\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4110__A1 _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5976__B _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5468__S _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5695__C _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5267__I _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4171__I _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5677__A1 _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5429__A1 _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6047__B _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_clk_i clknet_4_4_0_clk_i clknet_leaf_40_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6762__S _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_55_clk_i clknet_4_5_0_clk_i clknet_leaf_55_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4282__S _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5740_ memory\[23\]\[9\] _2247_ _2347_ _2205_ _2348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5671_ _1855_ _2257_ _2279_ _2280_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7410_ _3685_ _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_72_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4081__I net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8390_ _0690_ clknet_leaf_124_clk_i memory\[16\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4622_ memory\[22\]\[1\] _1173_ _1524_ _1526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_163_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7341_ _3660_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4553_ memory\[21\]\[1\] _1173_ _1487_ _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7272_ _1116_ memory\[3\]\[9\] _3614_ _3624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4484_ memory\[20\]\[1\] _1173_ _1450_ _1452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__I0 _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5668__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6223_ _2805_ _2810_ _2815_ _2820_ _2403_ _2821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_111_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6154_ _2529_ memory\[29\]\[18\] _2752_ _2389_ _2753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4340__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6085_ _2310_ memory\[11\]\[16\] _2685_ _2640_ _2686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5640__I _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5105_ _1242_ memory\[2\]\[1\] _1783_ _1785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4457__S _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5140__I0 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5036_ _1748_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5840__A1 _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_88_clk_i_I clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6987_ memory\[13\]\[3\] _1177_ _3469_ _3473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_137_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5938_ _2160_ memory\[19\]\[13\] _2540_ _2541_ _2542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4192__S _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8726_ _1026_ clknet_leaf_190_clk_i memory\[6\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_101_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8657_ _0957_ clknet_leaf_64_clk_i memory\[10\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5869_ _2467_ _2469_ _2471_ _2474_ _2475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__6148__A2 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7608_ _3802_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8588_ _0888_ clknet_leaf_91_clk_i memory\[4\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_2_0_clk_i clknet_0_clk_i clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7539_ memory\[5\]\[6\] net34 _3759_ _3766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_105_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4954__I0 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7008__S _3480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5659__A1 _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4706__I0 _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput45 net45 data_o[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_102_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput67 net67 data_o[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput56 net56 data_o[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__6847__S _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4367__S _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6084__A1 _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7120__I1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7678__S _3837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5831__A1 _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4166__I net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5198__S _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_119_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5198__I0 _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__S _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5898__A1 _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6330__B _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5725__I _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5661__S _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6757__S _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6075__A1 _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7890_ _0190_ clknet_leaf_74_clk_i memory\[18\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6910_ _3431_ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6841_ _1162_ memory\[9\]\[31\] _3360_ _3395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3984_ _1151_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6772_ _1954_ _3336_ _3356_ _3357_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_45_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8511_ _0811_ clknet_leaf_170_clk_i memory\[11\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5723_ _1855_ _2304_ _2329_ _2331_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__7178__I1 _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5654_ memory\[8\]\[7\] memory\[9\]\[7\] _1935_ _2264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5189__I0 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4740__S _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8442_ _0742_ clknet_leaf_217_clk_i memory\[13\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6240__B _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4605_ memory\[21\]\[26\] _1225_ _1509_ _1516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8373_ _0673_ clknet_leaf_187_clk_i memory\[14\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7324_ _1100_ memory\[4\]\[1\] _3650_ _3652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5585_ _1857_ _2192_ _2194_ _2195_ _2196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_130_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4536_ memory\[20\]\[26\] _1225_ _1472_ _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_68_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7255_ _3615_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4467_ _1080_ memory\[1\]\[26\] _1435_ _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6206_ _2803_ _2526_ memory\[25\]\[19\] _2804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5510__B1 _2117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7186_ _1093_ memory\[8\]\[0\] _3578_ _3579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4398_ _1080_ memory\[18\]\[26\] _1398_ _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6137_ memory\[2\]\[17\] memory\[3\]\[17\] _2736_ _2737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6066__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5113__I0 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7102__I1 _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6068_ memory\[22\]\[16\] _2669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5813__A1 _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5019_ memory\[27\]\[25\] _1223_ _1733_ _1739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8709_ _1009_ clknet_leaf_119_clk_i memory\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5973__C _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4927__I0 _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4097__S _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_111_clk_i_I clknet_4_15_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5280__I _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5804__A1 _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_17_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6907__I1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_36_clk_i_I clknet_4_4_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5370_ _1983_ _1985_ _1939_ _1986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_121_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4321_ _1362_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4252_ _1074_ memory\[29\]\[23\] _1322_ _1326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7040_ _3500_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_26_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6296__A1 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6219__C _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4183_ _1286_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7942_ _0242_ clknet_leaf_160_clk_i memory\[20\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6235__B _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7873_ _0173_ clknet_leaf_178_clk_i memory\[18\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6950__S _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6824_ _3386_ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_35_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3967_ _1097_ _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6755_ _1988_ memory\[10\]\[31\] _3341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_116_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5706_ memory\[8\]\[8\] memory\[9\]\[8\] _2314_ _2315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6771__A2 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3898_ _1091_ memory\[7\]\[31\] _1087_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6686_ _3258_ _3263_ _3268_ _3273_ _2894_ _3274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_8425_ _0725_ clknet_leaf_154_clk_i memory\[13\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5637_ _1895_ _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5326__A3 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7571__I1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5568_ _1988_ memory\[0\]\[5\] _2180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_14_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8356_ _0656_ clknet_leaf_158_clk_i memory\[14\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4519_ memory\[20\]\[18\] _1208_ _1461_ _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8287_ _0587_ clknet_leaf_180_clk_i memory\[30\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_44_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7307_ _3642_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5499_ _1883_ _2111_ _1887_ _2112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7238_ _1150_ memory\[8\]\[25\] _3600_ _3606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6039__A1 _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6129__C _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7169_ _3569_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4645__S _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5968__C _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_53_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6211__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5984__B _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7562__I1 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_5_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6039__C _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4619__I _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4555__S _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6825__I0 _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4870_ _1659_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7250__I0 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4290__S _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6540_ _3116_ _3121_ _3125_ _3130_ _2869_ _3131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6753__A2 _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6502__C _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6471_ memory\[4\]\[24\] _2934_ _3064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8210_ _0510_ clknet_leaf_33_clk_i memory\[28\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5422_ _1930_ memory\[10\]\[2\] _2037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_3_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8141_ _0441_ clknet_leaf_56_clk_i memory\[26\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5353_ memory\[23\]\[1\] _1896_ _1968_ _1899_ _1969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4304_ _1353_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7106__S _3528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8072_ _0372_ clknet_leaf_154_clk_i memory\[24\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5284_ _1058_ _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4235_ _1271_ memory\[29\]\[15\] _1311_ _1317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7023_ memory\[13\]\[20\] _1212_ _3491_ _3492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4166_ net15 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6816__I0 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4465__S _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6441__A1 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4097_ memory\[12\]\[28\] _1229_ _1213_ _1230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7925_ _0225_ clknet_leaf_195_clk_i memory\[1\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7856_ _0156_ clknet_leaf_71_clk_i memory\[17\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6807_ _3377_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4999_ _1728_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_108_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7787_ _0087_ clknet_leaf_77_clk_i memory\[15\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6744__A2 _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6738_ memory\[30\]\[31\] memory\[31\]\[31\] _1923_ _3324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6669_ memory\[15\]\[29\] _1896_ _3256_ _1899_ _3257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8408_ _0708_ clknet_leaf_24_clk_i memory\[16\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8339_ _0639_ clknet_leaf_80_clk_i memory\[9\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7016__S _3480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6855__S _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4530__I1 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4375__S _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6432__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7686__S _3837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7232__I0 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4597__I1 _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_209_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4521__I1 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6671__A1 _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4020_ memory\[12\]\[3\] _1177_ _1171_ _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5971_ _1863_ _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4922_ _1687_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8690_ _0990_ clknet_leaf_76_clk_i memory\[5\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4084__I net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7710_ _0010_ clknet_leaf_196_clk_i memory\[7\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7223__I0 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7641_ memory\[6\]\[22\] net20 _3817_ _3820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4853_ _1263_ memory\[25\]\[11\] _1649_ _1651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6726__A2 _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4784_ _1614_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4588__I1 _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6232__C _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7572_ _3783_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6523_ _2848_ memory\[27\]\[26\] _3113_ _2850_ _3114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_7_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6454_ _2629_ _3046_ _2961_ _3047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5405_ _1883_ _2019_ _1887_ _2020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6385_ memory\[4\]\[22\] _2934_ _2980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5336_ _1928_ _1940_ _1945_ _1951_ _1952_ _1953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_8124_ _0424_ clknet_leaf_7_clk_i memory\[25\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8055_ _0355_ clknet_leaf_41_clk_i memory\[23\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5267_ _1059_ _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7006_ memory\[13\]\[12\] _1196_ _3480_ _3483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_126_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4218_ _1254_ memory\[29\]\[7\] _1300_ _1308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6662__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5198_ _1125_ memory\[30\]\[13\] _1830_ _1834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input27_I data_i[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_5_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4149_ _1265_ memory\[15\]\[12\] _1261_ _1266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_158_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4276__I0 _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5311__C _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7462__I0 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4923__S _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7908_ _0208_ clknet_leaf_145_clk_i memory\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7839_ _0139_ clknet_leaf_182_clk_i memory\[29\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6423__B _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6142__C _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_210_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6653__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4503__I1 _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6317__C _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5929__S _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5392__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4990__I1 _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6170_ _2765_ _2767_ _2768_ _2769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5121_ _1258_ memory\[2\]\[9\] _1783_ _1793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6495__S _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7692__I0 _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3912__S _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5447__A2 _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_127_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5052_ _1756_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4003_ net6 _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_27_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4258__I0 _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7444__I0 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8742_ _1042_ clknet_leaf_107_clk_i memory\[7\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5954_ memory\[2\]\[13\] memory\[3\]\[13\] _2270_ _2558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5885_ memory\[23\]\[12\] _2247_ _2489_ _2205_ _2490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8673_ _0973_ clknet_leaf_146_clk_i memory\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4905_ _1678_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7624_ memory\[6\]\[14\] net11 _3806_ _3811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4836_ _1246_ memory\[25\]\[3\] _1638_ _1642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7555_ _3774_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6506_ _2779_ _3097_ _1994_ _3098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4767_ _1605_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7486_ _3737_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4698_ _1248_ memory\[23\]\[4\] _1562_ _1567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4981__I1 _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_84_clk_i_I clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6437_ memory\[24\]\[24\] _2799_ _3030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6368_ _2959_ _2962_ _2768_ _2963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8107_ _0407_ clknet_leaf_46_clk_i memory\[25\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5319_ memory\[8\]\[0\] memory\[9\]\[0\] _1935_ _1936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_54_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5438__A2 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6299_ _2796_ net51 _2896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6635__A1 _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8038_ _0338_ clknet_leaf_162_clk_i memory\[23\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4110__A2 _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4653__S _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5548__I _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4421__I0 _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7204__S _3578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4563__S _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5886__C _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5670_ _1954_ net68 _2280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4621_ _1525_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7340_ _1116_ memory\[4\]\[9\] _3650_ _3660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_52_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4552_ _1488_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7271_ _3623_ _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4483_ _1451_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6222_ _2817_ _2819_ _2768_ _2820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6153_ _2574_ memory\[28\]\[18\] _2752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4738__S _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7114__S _3505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6084_ _2362_ memory\[10\]\[16\] _2685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7665__I0 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6617__B2 _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5104_ _1784_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5035_ _1237_ memory\[28\]\[0\] _1747_ _1748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7417__I0 _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4473__S _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6986_ _3472_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5937_ _1866_ _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_0_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8725_ _1025_ clknet_leaf_188_clk_i memory\[6\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8656_ _0956_ clknet_leaf_65_clk_i memory\[10\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5868_ _2472_ _2473_ memory\[5\]\[11\] _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_7607_ memory\[6\]\[6\] net34 _3795_ _3802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_101_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_134_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8587_ _0887_ clknet_leaf_91_clk_i memory\[4\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5799_ _1893_ _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4819_ _1632_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5356__A1 _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7538_ _3765_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6420__C _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7469_ _3728_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput46 net46 data_o[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput57 net57 data_o[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput68 net68 data_o[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6608__A1 _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6863__S _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output58_I net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7408__I0 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4890__I0 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4383__S _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_184_clk_i clknet_4_3_0_clk_i clknet_leaf_184_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_27_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7694__S _3837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5278__I _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5595__B2 _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5347__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_199_clk_i clknet_4_2_0_clk_i clknet_leaf_199_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_91_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_122_clk_i clknet_4_14_0_clk_i clknet_leaf_122_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_137_clk_i clknet_4_9_0_clk_i clknet_leaf_137_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6870__I1 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_32_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4293__S _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6840_ _3394_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5586__A1 _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6771_ _1854_ net63 _3357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5722_ _2330_ net69 _2331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3983_ memory\[19\]\[25\] _1150_ _1140_ _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8510_ _0810_ clknet_leaf_169_clk_i memory\[11\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_99_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5653_ _1929_ memory\[11\]\[7\] _2262_ _2174_ _2263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5338__A1 _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8441_ _0741_ clknet_leaf_219_clk_i memory\[13\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8372_ _0672_ clknet_leaf_27_clk_i memory\[14\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4604_ _1515_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5584_ _1871_ _2060_ memory\[25\]\[6\] _2195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6948__S _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4535_ _1478_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7323_ _3651_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7254_ _1093_ memory\[3\]\[0\] _3614_ _3615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4466_ _1441_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7185_ _3577_ _3578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6205_ _1870_ _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_68_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5510__A1 _2107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4397_ _1404_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6136_ _1910_ _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6066__A2 _2665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6067_ _2664_ _2667_ _2291_ _2668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4872__I0 _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5018_ _1738_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6861__I1 _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5577__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4931__S _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6969_ _1154_ memory\[16\]\[27\] _3455_ _3463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_24_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8708_ _1008_ clknet_leaf_119_clk_i memory\[6\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5826__I _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5329__A1 _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8639_ _0939_ clknet_leaf_173_clk_i memory\[0\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6150__C _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5762__S _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_54_clk_i clknet_4_5_0_clk_i clknet_leaf_54_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_73_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6057__A2 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_69_clk_i clknet_4_7_0_clk_i clknet_leaf_69_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4863__I0 _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_125_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5568__A1 _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5002__S _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4091__I1 _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4640__I _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5740__B2 _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4320_ _1074_ memory\[17\]\[23\] _1358_ _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4288__S _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4251_ _1325_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I address_i[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7599__S _3795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4087__I net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4182_ _1078_ memory\[15\]\[25\] _1280_ _1286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7096__I1 _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7941_ _0241_ clknet_leaf_160_clk_i memory\[20\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7872_ _0172_ clknet_leaf_181_clk_i memory\[17\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6823_ _1144_ memory\[9\]\[22\] _3383_ _3386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5559__B2 _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4082__I1 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6754_ _3337_ _1894_ _3339_ _1901_ _3340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3966_ net18 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5705_ _1910_ _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6685_ _2933_ _3269_ _3271_ _3272_ _3273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_116_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4550__I _1486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7020__I1 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5636_ memory\[22\]\[7\] _2246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8424_ _0724_ clknet_leaf_150_clk_i memory\[13\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3897_ net30 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5567_ _2175_ _2178_ _1939_ _2179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5731__A1 _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6678__S _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8355_ _0655_ clknet_leaf_157_clk_i memory\[14\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4518_ _1469_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ memory\[30\]\[4\] memory\[31\]\[4\] _2066_ _2111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8286_ _0586_ clknet_leaf_189_clk_i memory\[30\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7306_ _1150_ memory\[3\]\[25\] _3636_ _3642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4449_ _1432_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5381__I _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7237_ _3605_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_129_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7168_ memory\[11\]\[24\] _1221_ _3564_ _3569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7087__I1 _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6119_ _2626_ memory\[19\]\[17\] _2718_ _2541_ _2719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7099_ _3532_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7302__S _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_12_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6145__C _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5757__S _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5970__A1 _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4073__I1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5722__A1 _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6278__A2 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_9_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_205_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5089__I0 _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4836__S _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5789__B2 _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6450__A2 _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4836__I0 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6336__B _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6202__A2 _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5961__A1 _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7002__I1 _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6470_ _3060_ _3062_ _2887_ _3063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_27_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5713__A1 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3915__S _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5421_ _2033_ _1921_ _2035_ _1927_ _2036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_40_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8140_ _0440_ clknet_leaf_55_clk_i memory\[26\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5352_ memory\[20\]\[1\] memory\[21\]\[1\] _1897_ _1968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4303_ _1271_ memory\[17\]\[15\] _1347_ _1353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5415__B _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6297__I _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8071_ _0371_ clknet_leaf_154_clk_i memory\[24\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5283_ memory\[23\]\[0\] _1896_ _1898_ _1899_ _1900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7022_ _3468_ _3491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4234_ _1316_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4165_ _1276_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4746__S _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7122__S _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6961__S _3455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4096_ net26 _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7924_ _0224_ clknet_leaf_81_clk_i memory\[1\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7855_ _0155_ clknet_leaf_89_clk_i memory\[17\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6806_ _1127_ memory\[9\]\[14\] _3372_ _3377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_34_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4998_ memory\[27\]\[15\] _1202_ _1722_ _1728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7786_ _0086_ clknet_leaf_178_clk_i memory\[15\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5952__A1 _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3949_ memory\[19\]\[14\] _1127_ _1119_ _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6737_ _2000_ memory\[29\]\[31\] _3322_ _1925_ _3323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5376__I _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6668_ memory\[12\]\[29\] memory\[13\]\[29\] _2919_ _3256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_1_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5619_ _2096_ memory\[6\]\[6\] _2230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8407_ _0707_ clknet_leaf_23_clk_i memory\[16\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_154_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6599_ _2981_ memory\[7\]\[27\] _3188_ _2983_ _3189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8338_ _0638_ clknet_leaf_95_clk_i memory\[9\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8269_ _0569_ clknet_leaf_61_clk_i memory\[30\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output40_I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6432__A2 _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_79_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5995__B _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7207__S _3589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6066__B _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ _2332_ _2569_ _2571_ _2572_ _2573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_99_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6781__S _3361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4921_ _1263_ memory\[26\]\[11\] _1685_ _1687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4852_ _1650_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6187__A1 _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7640_ _3819_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5934__B2 _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4783_ memory\[24\]\[10\] _1191_ _1613_ _1614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7571_ memory\[5\]\[21\] net19 _3781_ _3783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_99_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6522_ _2898_ memory\[26\]\[26\] _3113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_16_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6453_ memory\[16\]\[24\] memory\[17\]\[24\] _2630_ _3046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6021__S _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5404_ memory\[30\]\[2\] memory\[31\]\[2\] _1885_ _2019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8123_ _0423_ clknet_leaf_7_clk_i memory\[25\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6384_ _2976_ _2978_ _2887_ _2979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5335_ _1063_ _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8054_ _0354_ clknet_leaf_38_clk_i memory\[23\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5266_ _1882_ _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7005_ _3482_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4217_ _1307_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5870__B1 _2466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5197_ _1833_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4148_ net9 _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_97_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_80_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4079_ memory\[12\]\[22\] _1217_ _1213_ _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7907_ _0207_ clknet_leaf_145_clk_i memory\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6178__A1 _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7838_ _0138_ clknet_leaf_21_clk_i memory\[29\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5225__I0 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6973__I0 _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7769_ _0069_ clknet_leaf_219_clk_i memory\[12\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_137_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7027__S _3491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6350__A1 _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6866__S _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4386__S _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6614__B _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6333__C _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5392__A2 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6341__A1 _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5680__S _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5120_ _1792_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_71_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5051_ _1256_ memory\[28\]\[8\] _1747_ _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4002_ _1163_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_102_clk_i_I clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5412__C _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7400__S _3686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8741_ _1041_ clknet_leaf_117_clk_i memory\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5953_ _2267_ memory\[1\]\[13\] _2556_ _2509_ _2557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5884_ memory\[20\]\[12\] memory\[21\]\[12\] _2346_ _2489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6243__C _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_80_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8672_ _0972_ clknet_leaf_170_clk_i memory\[10\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4904_ _1246_ memory\[26\]\[3\] _1674_ _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5907__A1 _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7623_ _3810_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_103_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6955__I0 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4835_ _1641_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7554_ memory\[5\]\[13\] net10 _3770_ _3774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5383__A2 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ memory\[24\]\[2\] _1175_ _1602_ _1605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6580__A1 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6505_ memory\[8\]\[25\] memory\[9\]\[25\] _2780_ _3097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7485_ _1125_ memory\[10\]\[13\] _3733_ _3737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_27_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4697_ _1566_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6436_ _2846_ _3008_ _3028_ _3029_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6332__A1 _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7380__I0 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6367_ _2629_ _2960_ _2961_ _2962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4194__I0 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5318_ _1910_ _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_101_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8106_ _0406_ clknet_leaf_130_clk_i memory\[25\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_54_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6298_ _2875_ _2881_ _2888_ _2893_ _2894_ _2895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5249_ _1060_ _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8037_ _0337_ clknet_leaf_162_clk_i memory\[23\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6418__C _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6399__A1 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_119_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7310__S _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6946__I0 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5992__C _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6571__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_128_Left_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6328__C _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4488__I1 _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_137_Left_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4844__S _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6063__C _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4620_ memory\[22\]\[0\] _1164_ _1524_ _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5365__A2 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4551_ memory\[21\]\[0\] _1164_ _1487_ _1488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7270_ _1114_ memory\[3\]\[8\] _3614_ _3623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_80_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6314__B2 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4482_ memory\[20\]\[0\] _1164_ _1450_ _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6221_ _2629_ _2818_ _2495_ _2819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4176__I0 _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6152_ _2332_ _2747_ _2749_ _2750_ _2751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_57_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5103_ _1237_ memory\[2\]\[0\] _1783_ _1784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6083_ _2681_ _2406_ _2683_ _2360_ _2684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6617__A2 _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5034_ _1746_ _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4754__S _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7130__S _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6985_ memory\[13\]\[2\] _1175_ _3469_ _3472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5936_ _2208_ memory\[18\]\[13\] _2540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8724_ _1024_ clknet_leaf_79_clk_i memory\[6\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8655_ _0955_ clknet_leaf_94_clk_i memory\[10\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4651__I1 _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7606_ _3801_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5867_ _2006_ _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_8_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5798_ memory\[14\]\[10\] _2405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8586_ _0886_ clknet_leaf_87_clk_i memory\[4\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4818_ memory\[24\]\[27\] _1227_ _1624_ _1632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6553__A1 _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7537_ memory\[5\]\[5\] net33 _3759_ _3765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4749_ _1593_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5384__I _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7353__I0 _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7468_ _1108_ memory\[10\]\[5\] _3722_ _3728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6305__A1 _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4929__S _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4167__I0 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6419_ _2828_ memory\[10\]\[23\] _3013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_102_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput47 net47 data_o[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_7399_ _3691_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput58 net58 data_o[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput69 net69 data_o[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6608__A2 _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4664__S _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5595__A2 _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6919__I0 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6611__C _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5508__B _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5294__I _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4158__I0 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7215__S _3589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7647__I1 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4574__S _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__B2 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4330__I0 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5897__C _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3982_ net23 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6770_ _3340_ _3345_ _3350_ _3355_ _1063_ _3356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5721_ _1854_ _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_116_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3918__S _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5652_ _1930_ memory\[10\]\[7\] _2262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6535__A1 _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8440_ _0740_ clknet_leaf_218_clk_i memory\[13\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8371_ _0671_ clknet_leaf_78_clk_i memory\[14\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4603_ memory\[21\]\[25\] _1223_ _1509_ _1515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5583_ _1862_ memory\[27\]\[6\] _2193_ _1867_ _2194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_7322_ _1093_ memory\[4\]\[0\] _3650_ _3651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4534_ memory\[20\]\[25\] _1223_ _1472_ _1478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4149__I0 _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7253_ _3613_ _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4465_ _1078_ memory\[1\]\[25\] _1435_ _1441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6204_ _2382_ memory\[27\]\[19\] _2801_ _2384_ _2802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7184_ _1598_ _3359_ _3577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4396_ _1078_ memory\[18\]\[25\] _1398_ _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6135_ _2733_ memory\[1\]\[17\] _2734_ _2509_ _2735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6066_ _2288_ _2665_ _2666_ _2667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_84_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5017_ memory\[27\]\[24\] _1221_ _1733_ _1738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4484__S _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6774__A1 _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8707_ _1007_ clknet_leaf_144_clk_i memory\[6\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6968_ _3462_ _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4624__I1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5919_ memory\[24\]\[13\] _2333_ _2523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7594__I _3794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6899_ memory\[14\]\[26\] _1225_ _3419_ _3426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6526__A1 _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8638_ _0938_ clknet_leaf_171_clk_i memory\[0\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6431__C _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4388__I0 _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8569_ _0869_ clknet_leaf_204_clk_i memory\[3\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7326__I0 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4659__S _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7035__S _3491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output70_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6159__B _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6874__S _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4394__S _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_149_clk_i_I clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5510__C _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4615__I1 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6622__B _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6114__S _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6341__C _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_201_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6517__A1 _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4379__I0 _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5740__A2 _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4569__S _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5752__I _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4250_ _1072_ memory\[29\]\[22\] _1322_ _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4181_ _1285_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4303__I0 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7940_ _0240_ clknet_leaf_161_clk_i memory\[20\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7871_ _0171_ clknet_leaf_182_clk_i memory\[17\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6822_ _3385_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5559__A2 _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6756__A1 _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3965_ _1138_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6753_ memory\[15\]\[31\] _1896_ _3338_ _1899_ _3339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5704_ _1872_ _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6508__A1 _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6684_ _2938_ _2939_ memory\[5\]\[29\] _3272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3896_ _1090_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5635_ _2242_ _2244_ _1890_ _2245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6959__S _3455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8423_ _0723_ clknet_leaf_150_clk_i memory\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5031__I1 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5566_ _1934_ _2176_ _2177_ _2178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7308__I0 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8354_ _0654_ clknet_leaf_156_clk_i memory\[14\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4517_ memory\[20\]\[17\] _1206_ _1461_ _1469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5497_ _2063_ memory\[29\]\[4\] _2109_ _1880_ _2110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7305_ _3641_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8285_ _0585_ clknet_leaf_190_clk_i memory\[30\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4448_ _1275_ memory\[1\]\[17\] _1424_ _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7236_ _1148_ memory\[8\]\[24\] _3600_ _3605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_183_clk_i clknet_4_3_0_clk_i clknet_leaf_183_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_0_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_129_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4379_ _1275_ memory\[18\]\[17\] _1387_ _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7167_ _3568_ _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6118_ _2674_ memory\[18\]\[17\] _2718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6707__B _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7098_ memory\[31\]\[23\] _1219_ _3528_ _3532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6049_ memory\[4\]\[15\] _2468_ _2651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5611__B _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5103__S _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_198_clk_i clknet_4_2_0_clk_i clknet_leaf_198_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_150_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5330__C _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4942__S _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_121_clk_i clknet_4_11_0_clk_i clknet_leaf_121_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_37_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_136_clk_i clknet_4_9_0_clk_i clknet_leaf_136_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_134_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__A2 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_75_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5486__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7499__I _3721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5789__A2 _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6109__S _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5013__S _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__A2 _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5013__I1 _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6779__S _3361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5420_ memory\[15\]\[2\] _1922_ _2034_ _1925_ _2035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4299__S _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5482__I _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5351_ memory\[22\]\[1\] _1967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4302_ _1352_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8070_ _0370_ clknet_leaf_156_clk_i memory\[24\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5282_ _1879_ _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4233_ _1269_ memory\[29\]\[14\] _1311_ _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7021_ _3490_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_57_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__A1 _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4164_ _1275_ memory\[15\]\[17\] _1261_ _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_65_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4095_ _1228_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5431__B _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7923_ _0223_ clknet_leaf_83_clk_i memory\[1\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6246__C _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5858__S _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7854_ _0154_ clknet_leaf_101_clk_i memory\[17\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6729__A1 _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4762__S _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6805_ _3376_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5657__I _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6262__B _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7785_ _0085_ clknet_leaf_153_clk_i memory\[15\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_53_clk_i clknet_4_5_0_clk_i clknet_leaf_53_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4997_ _1727_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6736_ _2001_ memory\[28\]\[31\] _3322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5401__A1 _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3948_ net11 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5004__I1 _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5593__S _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3879_ _1078_ memory\[7\]\[25\] _1066_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6667_ memory\[14\]\[29\] _3255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5618_ memory\[4\]\[6\] _1998_ _2229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8406_ _0706_ clknet_leaf_25_clk_i memory\[16\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6598_ _1864_ memory\[6\]\[27\] _3188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8337_ _0637_ clknet_leaf_96_clk_i memory\[9\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_68_clk_i clknet_4_13_0_clk_i clknet_leaf_68_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5549_ _1905_ memory\[18\]\[5\] _2161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_42_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3905__I _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8268_ _0568_ clknet_leaf_58_clk_i memory\[30\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7219_ _1131_ memory\[8\]\[16\] _3589_ _3596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4937__S _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8199_ _0499_ clknet_leaf_128_clk_i memory\[28\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_100_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4818__I1 _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4672__S _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6991__I1 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4754__I0 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7223__S _3589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7022__I _3468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5631__A1 _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4582__S _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4920_ _1686_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4851_ _1260_ memory\[25\]\[10\] _1649_ _1650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_136_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5934__A2 _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4782_ _1601_ _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7570_ _3782_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_99_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ memory\[24\]\[26\] _2799_ _3112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6452_ _2626_ memory\[19\]\[24\] _3044_ _2003_ _3045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5403_ _1876_ memory\[29\]\[2\] _2017_ _1880_ _2018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5426__B _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8122_ _0422_ clknet_leaf_7_clk_i memory\[25\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6383_ _2884_ _2977_ _2602_ _2978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5334_ _1947_ _1949_ _1950_ _1951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5265_ _1060_ _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8053_ _0353_ clknet_leaf_36_clk_i memory\[23\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7004_ memory\[13\]\[11\] _1194_ _3480_ _3482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5196_ _1123_ memory\[30\]\[12\] _1830_ _1833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4216_ _1252_ memory\[29\]\[6\] _1300_ _1307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4147_ _1264_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5622__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5588__S _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_23_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4078_ net20 _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_108_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7906_ _0206_ clknet_leaf_141_clk_i memory\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4492__S _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7837_ _0137_ clknet_leaf_16_clk_i memory\[29\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6704__C _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5387__I _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7768_ _0068_ clknet_leaf_218_clk_i memory\[12\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_137_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7699_ _3849_ _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6719_ _1904_ memory\[1\]\[30\] _3305_ _2975_ _3306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_117_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7308__S _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5689__A1 _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4736__I0 _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6102__A2 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5161__I0 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7043__S _3468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6882__S _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5498__S _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5613__A1 _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4727__I0 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7141__I1 _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5050_ _1755_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5852__A1 _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6077__B _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4001_ memory\[19\]\[31\] _1162_ _1097_ _1163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5952_ _2318_ memory\[0\]\[13\] _2556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_88_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8740_ _1040_ clknet_leaf_118_clk_i memory\[7\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_197_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4903_ _1677_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5883_ memory\[22\]\[12\] _2488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8671_ _0971_ clknet_leaf_170_clk_i memory\[10\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7622_ memory\[6\]\[13\] net10 _3806_ _3810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4834_ _1244_ memory\[25\]\[2\] _1638_ _1641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7553_ _3773_ _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_103_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4765_ _1604_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7128__S _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ _2776_ memory\[11\]\[25\] _3095_ _1907_ _3096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_7484_ _3736_ _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4696_ _1246_ memory\[23\]\[3\] _1562_ _1566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6967__S _3455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6435_ _2796_ net54 _3029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_132_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6366_ _1057_ _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5317_ _1872_ _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_54_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8105_ _0405_ clknet_leaf_177_clk_i memory\[25\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7132__I1 _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6096__A1 _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8036_ _0336_ clknet_leaf_161_clk_i memory\[23\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6297_ _1063_ _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5843__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input32_I data_i[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5603__C _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5248_ _1864_ memory\[26\]\[0\] _1865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5179_ _1106_ memory\[30\]\[4\] _1819_ _1824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5111__S _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6434__C _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4950__S _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5134__I0 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6087__A1 _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5834__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4196__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5021__S _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6011__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__I0 _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4550_ _1486_ _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_13_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6787__S _3361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5691__S _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6314__A2 _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4481_ _1449_ _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_13_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6220_ memory\[16\]\[19\] memory\[17\]\[19\] _2630_ _2818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6151_ _2337_ _2526_ memory\[25\]\[18\] _2750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5102_ _1782_ _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7114__I1 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4100__S _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6082_ memory\[15\]\[16\] _2357_ _2682_ _2307_ _2683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5423__C _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5033_ _1598_ _1294_ _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__7411__S _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6254__C _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6984_ _3471_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5935_ _2536_ _2294_ _2538_ _2250_ _2539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8723_ _1023_ clknet_leaf_78_clk_i memory\[6\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4100__I1 _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8654_ _0954_ clknet_leaf_95_clk_i memory\[10\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5866_ _1870_ _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_8_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4770__S _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7605_ memory\[6\]\[5\] net33 _3795_ _3801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4817_ _1631_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8585_ _0885_ clknet_leaf_110_clk_i memory\[4\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5797_ _2387_ _2393_ _2397_ _2402_ _2403_ _2404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_90_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6270__B _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7536_ _3764_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4748_ _1084_ memory\[23\]\[28\] _1584_ _1593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4679_ _1555_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6305__A2 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7467_ _3727_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6418_ _3009_ _2872_ _3011_ _2826_ _3012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_113_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput48 net48 data_o[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7398_ _1106_ memory\[0\]\[4\] _3686_ _3691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6349_ memory\[24\]\[22\] _2799_ _2944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput59 net59 data_o[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_12_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8019_ _0319_ clknet_leaf_34_clk_i memory\[22\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_67_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6445__B _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6164__C _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4680__S _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6544__A2 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_145_clk_i_I clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5524__B _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5107__I0 _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4855__S _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5283__A2 _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6480__A1 _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6232__A1 _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3981_ _1149_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5720_ _2309_ _2317_ _2323_ _2328_ _1952_ _2329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__4590__S _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5686__S _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5651_ _2258_ _1921_ _2260_ _1927_ _2261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_26_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7583__I1 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8370_ _0670_ clknet_leaf_76_clk_i memory\[14\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4602_ _1514_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5582_ _1957_ memory\[26\]\[6\] _2193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7321_ _3649_ _3650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_81_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _1477_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7406__S _3686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7252_ _1062_ _1411_ _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__6299__A1 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6203_ _2432_ memory\[26\]\[19\] _2801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_68_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4464_ _1440_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4829__I _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4395_ _1403_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7183_ _3576_ _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6134_ _2318_ memory\[0\]\[17\] _2734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_111_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _1293_ _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7141__S _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5016_ _1737_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6967_ _1152_ memory\[16\]\[26\] _3455_ _3462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5918_ _2380_ _2498_ _2521_ _2522_ _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_8706_ _1006_ clknet_leaf_144_clk_i memory\[6\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6898_ _3425_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6712__C _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5849_ memory\[15\]\[11\] _2357_ _2454_ _2307_ _2455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_119_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8637_ _0937_ clknet_leaf_171_clk_i memory\[0\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_133_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8568_ _0868_ clknet_leaf_204_clk_i memory\[3\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7519_ _3754_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6220__S _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8499_ _0799_ clknet_leaf_78_clk_i memory\[11\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7316__S _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output63_I net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6954__I _3432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6837__I0 _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6462__A1 _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_71_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7262__I0 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6765__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__B _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6130__S _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4551__I1 _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4180_ _1076_ memory\[15\]\[24\] _1280_ _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7870_ _0170_ clknet_leaf_186_clk_i memory\[17\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6821_ _1142_ memory\[9\]\[21\] _3383_ _3385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3964_ memory\[19\]\[19\] _1137_ _1119_ _1138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6752_ memory\[12\]\[31\] memory\[13\]\[31\] _1897_ _3338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7556__I1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5703_ _2310_ memory\[11\]\[8\] _2311_ _2174_ _2312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_57_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6683_ _2981_ memory\[7\]\[29\] _3270_ _2983_ _3271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3895_ _1089_ memory\[7\]\[30\] _1087_ _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5634_ _1883_ _2243_ _2200_ _2244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8422_ _0722_ clknet_leaf_159_clk_i memory\[13\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8353_ _0653_ clknet_leaf_151_clk_i memory\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6040__S _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7136__S _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5565_ _1238_ _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5731__A3 _2336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7304_ _1148_ memory\[3\]\[24\] _3636_ _3641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4516_ _1468_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5496_ _2108_ memory\[28\]\[4\] _2109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8284_ _0584_ clknet_leaf_17_clk_i memory\[30\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4447_ _1431_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6975__S _3432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7235_ _3604_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4542__I1 _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6692__A1 _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7166_ memory\[11\]\[23\] _1219_ _3564_ _3568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_129_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4378_ _1394_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6117_ _2712_ _2294_ _2715_ _2716_ _2717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6819__I0 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7097_ _3531_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_13_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6048_ _2647_ _2649_ _2421_ _2650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_68_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7244__I0 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7999_ _0299_ clknet_leaf_81_clk_i memory\[21\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_37_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__S _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4758__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_18_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6683__A1 _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6435__A1 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7483__I0 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4297__I0 _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5521__C _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6633__B _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6125__S _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5410__A2 _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5350_ _1963_ _1965_ _1890_ _1966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__I1 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4301_ _1269_ memory\[17\]\[14\] _1347_ _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6795__S _3361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5281_ memory\[20\]\[0\] memory\[21\]\[0\] _1897_ _1898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4232_ _1315_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7020_ memory\[13\]\[19\] _1210_ _3480_ _3490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6674__A1 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4524__I1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5204__S _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4163_ net14 _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4288__I0 _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7474__I0 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6527__C _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4094_ memory\[12\]\[27\] _1227_ _1213_ _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7922_ _0222_ clknet_leaf_83_clk_i memory\[1\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7853_ _0153_ clknet_leaf_99_clk_i memory\[17\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6729__A2 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6804_ _1125_ memory\[9\]\[13\] _3372_ _3376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4996_ memory\[27\]\[14\] _1200_ _1722_ _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7784_ _0084_ clknet_leaf_151_clk_i memory\[15\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3947_ _1126_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6735_ _1887_ _3317_ _3319_ _3320_ _3321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_19_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6666_ _3239_ _3244_ _3248_ _3253_ _2869_ _3254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_46_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3878_ net23 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_116_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5617_ _2225_ _2227_ _1950_ _2228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4212__I0 _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8405_ _0705_ clknet_leaf_26_clk_i memory\[16\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6597_ memory\[4\]\[27\] _2934_ _3187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8336_ _0636_ clknet_leaf_96_clk_i memory\[9\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5548_ _1903_ _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_42_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8267_ _0567_ clknet_leaf_74_clk_i memory\[30\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7218_ _3595_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5479_ _1941_ _2092_ _1994_ _2093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4515__I1 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8198_ _0498_ clknet_leaf_128_clk_i memory\[28\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7149_ memory\[11\]\[15\] _1202_ _3553_ _3559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_70_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6417__B2 _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7217__I0 _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5784__S _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5516__C _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5459__A2 _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7504__S _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5251__C _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4863__S _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4690__I0 _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4850_ _1637_ _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_47_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_182_clk_i clknet_4_9_0_clk_i clknet_leaf_182_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5395__A1 _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4442__I0 _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4781_ _1612_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6520_ _2846_ _3090_ _3110_ _3111_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_7_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5707__B _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6451_ _2674_ memory\[18\]\[24\] _3044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_15_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5402_ _1877_ memory\[28\]\[2\] _2017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_42_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6382_ memory\[2\]\[22\] memory\[3\]\[22\] _2736_ _2977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4103__S _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_197_clk_i clknet_4_2_0_clk_i clknet_leaf_197_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_193_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5333_ _1915_ _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8121_ _0421_ clknet_leaf_9_clk_i memory\[25\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8052_ _0352_ clknet_leaf_34_clk_i memory\[23\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_120_clk_i clknet_4_14_0_clk_i clknet_leaf_120_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5264_ _1876_ memory\[29\]\[0\] _1878_ _1880_ _1881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6538__B _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5195_ _1832_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7003_ _3481_ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4215_ _1306_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4146_ _1263_ memory\[15\]\[11\] _1261_ _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_135_clk_i clknet_4_9_0_clk_i clknet_leaf_135_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_39_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4077_ _1216_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7905_ _0205_ clknet_leaf_140_clk_i memory\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7836_ _0136_ clknet_leaf_16_clk_i memory\[29\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5386__A1 _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4979_ memory\[27\]\[6\] _1183_ _1711_ _1718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7767_ _0067_ clknet_leaf_5_clk_i memory\[12\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_137_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7698_ _1135_ memory\[7\]\[18\] _1065_ _3849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6718_ _1905_ memory\[0\]\[30\] _3305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5617__B _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6649_ _2848_ memory\[27\]\[29\] _3236_ _2850_ _3237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_18_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5109__S _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5336__C _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7324__S _3650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8319_ _0619_ clknet_leaf_180_clk_i net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4948__S _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7686__I0 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7438__I0 _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6183__B _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6630__C _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4975__I1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5019__S _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7234__S _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6358__B _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6629__A1 _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_52_clk_i clknet_4_5_0_clk_i clknet_leaf_52_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7429__I0 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4000_ net30 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4593__S _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6093__B _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5951_ _2552_ _2554_ _2414_ _2555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_99_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_67_clk_i clknet_4_7_0_clk_i clknet_leaf_67_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8670_ _0970_ clknet_leaf_169_clk_i memory\[10\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4902_ _1244_ memory\[26\]\[2\] _1674_ _1677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5882_ _2484_ _2486_ _2291_ _2487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7621_ _3809_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3937__S _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4415__I0 _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4833_ _1640_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7552_ memory\[5\]\[12\] net9 _3770_ _3773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_103_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6313__S _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4764_ memory\[24\]\[1\] _1173_ _1602_ _1604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7483_ _1123_ memory\[10\]\[12\] _3733_ _3736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6540__C _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6503_ _2828_ memory\[10\]\[25\] _3095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4695_ _1565_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6434_ _3012_ _3017_ _3022_ _3027_ _2894_ _3028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_113_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5540__A1 _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6365_ memory\[16\]\[22\] memory\[17\]\[22\] _2630_ _2960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4768__S _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5316_ _1929_ memory\[11\]\[0\] _1931_ _1932_ _1933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6296_ _2467_ _2889_ _2891_ _2892_ _2893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_8104_ _0404_ clknet_leaf_138_clk_i memory\[25\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5247_ _1863_ _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6983__S _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8035_ _0335_ clknet_leaf_166_clk_i memory\[23\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5178_ _1823_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6891__I1 _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input25_I data_i[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4129_ net34 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_79_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7819_ _0119_ clknet_leaf_73_clk_i memory\[29\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4406__I0 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6450__C _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5531__A1 _2127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4678__S _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7054__S _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5861__I _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6893__S _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6882__I1 _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_141_clk_i_I clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5598__A1 _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5070__I0 _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6562__A3 _3151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5770__A1 _2361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4480_ _1169_ _1448_ _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_12_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_66_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4588__S _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6150_ _2382_ memory\[27\]\[18\] _2748_ _2384_ _2749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_21_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6088__B _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5101_ _1374_ _1411_ _1782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6081_ memory\[12\]\[16\] memory\[13\]\[16\] _2453_ _2682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5825__A2 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5032_ _1745_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4884__I0 _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6250__A2 _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6983_ memory\[13\]\[1\] _1173_ _3469_ _3471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5934_ memory\[23\]\[13\] _2247_ _2537_ _2205_ _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8722_ _1022_ clknet_leaf_76_clk_i memory\[6\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8653_ _0953_ clknet_leaf_95_clk_i memory\[10\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5865_ _2049_ memory\[7\]\[11\] _2470_ _2051_ _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_8_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6002__A2 _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7139__S _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4850__I _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7604_ _3800_ _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7050__I1 _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4816_ memory\[24\]\[26\] _1225_ _1624_ _1631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8584_ _0884_ clknet_leaf_107_clk_i memory\[4\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5796_ _1094_ _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5761__A1 _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7535_ memory\[5\]\[4\] net32 _3759_ _3764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4747_ _1592_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4678_ memory\[22\]\[28\] _1229_ _1546_ _1555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7466_ _1106_ memory\[10\]\[4\] _3722_ _3727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_116_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4498__S _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7397_ _3690_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5513__B2 _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6417_ memory\[15\]\[23\] _2823_ _3010_ _2773_ _3011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5614__C _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput49 net49 data_o[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6348_ _2846_ _2917_ _2942_ _2943_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_101_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6279_ _2828_ memory\[10\]\[20\] _2876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5816__A2 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8018_ _0318_ clknet_leaf_45_clk_i memory\[22\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_67_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6241__A2 _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7041__I1 _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7512__S _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_7_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6855__I1 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4000__I net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6355__C _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3980_ memory\[19\]\[24\] _1148_ _1140_ _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4094__I1 _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5991__A1 _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5650_ memory\[15\]\[7\] _1922_ _2259_ _1925_ _2260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__6090__C _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_100_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4601_ memory\[21\]\[24\] _1221_ _1509_ _1514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5043__I0 _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6791__I0 _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6798__S _3372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5743__A1 _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5581_ memory\[24\]\[6\] _1859_ _2192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4532_ memory\[20\]\[24\] _1221_ _1472_ _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7320_ _1238_ _1064_ _1598_ _3649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XPHY_EDGE_ROW_68_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6299__A2 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7251_ _3612_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4463_ _1076_ memory\[1\]\[24\] _1435_ _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6202_ memory\[24\]\[19\] _2799_ _2800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4394_ _1076_ memory\[18\]\[24\] _1398_ _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7182_ memory\[11\]\[31\] _1235_ _3541_ _3576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_68_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6133_ _1903_ _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6064_ memory\[30\]\[16\] memory\[31\]\[16\] _2532_ _2665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_111_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__I0 _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5015_ memory\[27\]\[23\] _1219_ _1733_ _1737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6471__A2 _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_77_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6966_ _3461_ _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5917_ _2330_ net42 _2522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8705_ _1005_ clknet_leaf_145_clk_i memory\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_24_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4085__I1 _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5982__A1 _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6897_ memory\[14\]\[25\] _1223_ _3419_ _3425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7023__I1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5848_ memory\[12\]\[11\] memory\[13\]\[11\] _2453_ _2454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5609__C _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8636_ _0936_ clknet_leaf_197_clk_i memory\[0\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5779_ _2337_ _2060_ memory\[25\]\[10\] _2386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_86_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8567_ _0867_ clknet_leaf_203_clk_i memory\[3\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7518_ _1158_ memory\[10\]\[29\] _3744_ _3754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8498_ _0798_ clknet_leaf_66_clk_i memory\[11\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5117__S _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7449_ _3717_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4956__S _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7332__S _3650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_95_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4848__I0 _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output56_I net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_14_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_129_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4076__I1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7014__I1 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A1 _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6411__S _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_136_Right_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5027__S _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6150__A1 _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7242__S _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6085__C _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6820_ _3384_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5697__S _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5964__A1 _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3963_ net16 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_46_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6751_ memory\[14\]\[31\] _3337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_116_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5702_ _1930_ memory\[10\]\[8\] _2311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_85_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5429__C _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3894_ net29 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4106__S _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6682_ _1864_ memory\[6\]\[29\] _3270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5716__A1 _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5633_ memory\[30\]\[7\] memory\[31\]\[7\] _2066_ _2243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8421_ _0721_ clknet_leaf_159_clk_i memory\[13\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7417__S _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5564_ memory\[8\]\[5\] memory\[9\]\[5\] _1935_ _2176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8352_ _0652_ clknet_leaf_167_clk_i memory\[9\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4515_ memory\[20\]\[16\] _1204_ _1461_ _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7303_ _3640_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5495_ _1863_ _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_14_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8283_ _0583_ clknet_leaf_3_clk_i memory\[30\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4446_ _1273_ memory\[1\]\[16\] _1424_ _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_113_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6141__A1 _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7234_ _1146_ memory\[8\]\[23\] _3600_ _3604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4377_ _1273_ memory\[18\]\[16\] _1387_ _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6692__A2 _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7165_ _3567_ _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4776__S _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _1058_ _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_119_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7096_ memory\[31\]\[22\] _1217_ _3528_ _3531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6047_ _2418_ _2648_ _2602_ _2649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6991__S _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_188_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7998_ _0298_ clknet_leaf_30_clk_i memory\[21\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5955__A1 _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6949_ _3452_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8619_ _0919_ clknet_leaf_104_clk_i memory\[0\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5707__A1 _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7062__S _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5802__C _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6435__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6199__A1 _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6406__S _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6205__I _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4300_ _1351_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5280_ _1884_ _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_121_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4231_ _1267_ memory\[29\]\[13\] _1311_ _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4162_ _1274_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4093_ net25 _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7921_ _0221_ clknet_leaf_90_clk_i memory\[1\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7852_ _0152_ clknet_leaf_103_clk_i memory\[17\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6803_ _3375_ _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4995_ _1726_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7783_ _0083_ clknet_leaf_151_clk_i memory\[15\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3946_ memory\[19\]\[13\] _1125_ _1119_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6734_ _1870_ _1990_ memory\[25\]\[31\] _3320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_34_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7147__S _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8404_ _0704_ clknet_leaf_28_clk_i memory\[16\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6665_ _3250_ _3252_ _1915_ _3253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_6_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3877_ _1077_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5616_ _1941_ _2226_ _2136_ _2227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6596_ _3183_ _3185_ _2887_ _3186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8335_ _0635_ clknet_leaf_97_clk_i memory\[9\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5547_ _2156_ _1894_ _2158_ _1901_ _2159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_8266_ _0566_ clknet_leaf_86_clk_i memory\[30\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5478_ memory\[2\]\[3\] memory\[3\]\[3\] _1992_ _2092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7217_ _1129_ memory\[8\]\[15\] _3589_ _3595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4429_ _1256_ memory\[1\]\[8\] _1413_ _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_57_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8197_ _0497_ clknet_leaf_129_clk_i memory\[28\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7148_ _3558_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7079_ memory\[31\]\[14\] _1200_ _3517_ _3522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6417__A2 _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5130__S _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6226__S _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6353__A1 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6105__A1 _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5813__B _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6628__C _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6408__A2 _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7520__S _3721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5219__I0 _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6967__I0 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4780_ memory\[24\]\[9\] _1189_ _1602_ _1612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6592__A1 _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6450_ _3040_ _2760_ _3042_ _2716_ _3043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7392__I0 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6344__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_136_clk_i_I clknet_4_9_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_41_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5401_ _1857_ _2012_ _2014_ _2015_ _2016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6381_ _2733_ memory\[1\]\[22\] _2974_ _2975_ _2976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5332_ _1934_ _1948_ _1887_ _1949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8120_ _0420_ clknet_leaf_9_clk_i memory\[25\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8051_ _0351_ clknet_leaf_42_clk_i memory\[23\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5263_ _1879_ _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_76_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5215__S _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6647__A2 _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5194_ _1121_ memory\[30\]\[11\] _1830_ _1832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7002_ memory\[13\]\[10\] _1191_ _3480_ _3481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4214_ _1250_ memory\[29\]\[5\] _1300_ _1306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4145_ net8 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_39_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6554__B _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4130__I0 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4076_ memory\[12\]\[21\] _1215_ _1213_ _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6046__S _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6273__C _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7904_ _0204_ clknet_leaf_134_clk_i memory\[18\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7835_ _0135_ clknet_leaf_16_clk_i memory\[29\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_121_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4978_ _1717_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7766_ _0066_ clknet_leaf_5_clk_i memory\[12\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_137_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3929_ net36 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7697_ _3848_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6717_ _3301_ _3303_ _1890_ _3304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_117_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6648_ _2898_ memory\[26\]\[29\] _3236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_6_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6335__A1 _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__S _3795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6579_ memory\[16\]\[27\] memory\[17\]\[27\] _1885_ _3169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8318_ _0618_ clknet_leaf_190_clk_i net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3932__I net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8249_ _0549_ clknet_leaf_204_clk_i memory\[2\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7340__S _3650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6464__B _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4121__I0 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4672__I1 _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5808__B _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5594__I _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4204__S _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7374__I0 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4188__I0 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5543__B _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5035__S _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4360__I0 _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__S _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7250__S _3577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5950_ _2313_ _2553_ _2177_ _2554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_62_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4112__I0 _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4901_ _1676_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5881_ _2288_ _2485_ _2200_ _2486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7620_ memory\[6\]\[12\] net9 _3806_ _3809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_62_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4832_ _1242_ memory\[25\]\[1\] _1638_ _1640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6565__A1 _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7551_ _3772_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_103_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4763_ _1603_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7482_ _3735_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5437__C _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6317__A1 _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4694_ _1244_ memory\[23\]\[2\] _1562_ _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6502_ _3091_ _2872_ _3093_ _2826_ _3094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_113_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6433_ _2933_ _3023_ _3025_ _3026_ _3027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_125_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7425__S _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6364_ _2626_ memory\[19\]\[22\] _2958_ _2541_ _2959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6549__B _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5315_ _1866_ _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6295_ _2472_ _2473_ memory\[5\]\[20\] _2892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8103_ _0403_ clknet_leaf_176_clk_i memory\[25\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5246_ _1059_ _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6268__C _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8034_ _0334_ clknet_leaf_165_clk_i memory\[23\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5177_ _1104_ memory\[30\]\[3\] _1819_ _1823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7160__S _3564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5679__I _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6284__B _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4128_ _1251_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4059_ net13 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_79_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input18_I data_i[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7818_ _0118_ clknet_leaf_82_clk_i memory\[29\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_65_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6556__A1 _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7749_ _0049_ clknet_leaf_159_clk_i memory\[12\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5347__C _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6308__A1 _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7659__I1 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_181_clk_i clknet_4_9_0_clk_i clknet_leaf_181_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4694__S _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5810__C _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5589__I _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4645__I1 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_196_clk_i clknet_4_2_0_clk_i clknet_leaf_196_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_84_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4270__A2 _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_106_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6641__C _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7347__I0 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4869__S _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_134_clk_i clknet_4_9_0_clk_i clknet_leaf_134_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_41_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_115_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6080_ memory\[14\]\[16\] _2681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5100_ _1781_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_57_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5031_ memory\[27\]\[31\] _1235_ _1710_ _1745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_149_clk_i clknet_4_11_0_clk_i clknet_leaf_149_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__C _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8721_ _1021_ clknet_leaf_69_clk_i memory\[6\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4636__I1 _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6982_ _3470_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5933_ memory\[20\]\[13\] memory\[21\]\[13\] _2346_ _2537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_124_Left_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8652_ _0952_ clknet_leaf_95_clk_i memory\[10\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5864_ _2096_ memory\[6\]\[11\] _2470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_91_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6551__C _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6324__S _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6538__A1 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8583_ _0883_ clknet_leaf_107_clk_i memory\[4\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7603_ memory\[6\]\[4\] net32 _3795_ _3800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4815_ _1630_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5795_ _2399_ _2401_ _2302_ _2402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_90_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7534_ _3763_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7338__I0 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4746_ _1082_ memory\[23\]\[27\] _1584_ _1592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7155__S _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4677_ _1554_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7465_ _3726_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_133_Left_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7396_ _1104_ memory\[0\]\[3\] _3686_ _3690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5513__A2 _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6416_ memory\[12\]\[23\] memory\[13\]\[23\] _2919_ _3010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput39 net39 data_o[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6347_ _2796_ net52 _2943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7510__I0 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6278_ _2871_ _2872_ _2874_ _2826_ _2875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8017_ _0317_ clknet_leaf_54_clk_i memory\[22\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4324__I0 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5229_ _1156_ memory\[30\]\[28\] _1841_ _1850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_67_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6529__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5358__B _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_51_clk_i clknet_4_5_0_clk_i clknet_leaf_51_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_124_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_10_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5504__A2 _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_66_clk_i clknet_4_7_0_clk_i clknet_leaf_66_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6189__B _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6701__B2 _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5540__C _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6768__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5440__A1 _2036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5983__S _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4600_ _1513_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_19_clk_i clknet_4_3_0_clk_i clknet_leaf_19_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_81_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5580_ _1855_ _2168_ _2190_ _2191_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_53_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5782__I _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4599__S _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4531_ _1476_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7250_ _1162_ memory\[8\]\[31\] _3577_ _3612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4462_ _1439_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6201_ _1858_ _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4393_ _1402_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7181_ _3575_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6132_ _2729_ _2731_ _2414_ _2732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_110_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6063_ _2529_ memory\[29\]\[16\] _2663_ _2389_ _2664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_84_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6456__B1 _3043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ _1736_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6546__C _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5223__S _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4609__I1 _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6965_ _1150_ memory\[16\]\[25\] _3455_ _3461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5431__A1 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5916_ _2502_ _2507_ _2513_ _2520_ _2428_ _2521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_24_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8704_ _1004_ clknet_leaf_179_clk_i memory\[5\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8635_ _0935_ clknet_leaf_207_clk_i memory\[0\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6896_ _3424_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_134_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7184__A1 _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5847_ _1884_ _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6989__S _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5778_ _2382_ memory\[27\]\[10\] _2383_ _2384_ _2385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8566_ _0866_ clknet_leaf_202_clk_i memory\[3\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8497_ _0797_ clknet_leaf_66_clk_i memory\[11\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4729_ _1056_ memory\[23\]\[19\] _1573_ _1583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7517_ _3753_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_184_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7448_ _1156_ memory\[0\]\[28\] _3708_ _3717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7613__S _3795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7379_ _3680_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_73_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__C _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5360__C _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output49_I net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5670__A1 _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6028__I _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5867__I _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5422__A1 _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6899__S _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5025__I1 _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4212__S _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5489__A1 _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3850__I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5043__S _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5978__S _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4882__S _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5777__I _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6750_ _3321_ _3326_ _3330_ _3335_ _1094_ _3336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5701_ _1903_ _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3962_ _1136_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6681_ memory\[4\]\[29\] _2934_ _3269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3893_ _1088_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5632_ _2063_ memory\[29\]\[7\] _2241_ _1880_ _2242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_72_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8420_ _0720_ clknet_leaf_158_clk_i memory\[13\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5563_ _1929_ memory\[11\]\[5\] _2173_ _2174_ _2175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8351_ _0651_ clknet_leaf_170_clk_i memory\[9\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4514_ _1467_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7302_ _1146_ memory\[3\]\[23\] _3636_ _3640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5445__C _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5494_ _1857_ _2103_ _2105_ _2106_ _2107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_8282_ _0582_ clknet_leaf_2_clk_i memory\[30\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4445_ _1430_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_113_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3961__S _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7233_ _3603_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4376_ _1393_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7164_ memory\[11\]\[22\] _1217_ _3564_ _3567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_129_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6115_ memory\[23\]\[17\] _2713_ _2714_ _2671_ _2715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7095_ _3530_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6046_ memory\[2\]\[15\] memory\[3\]\[15\] _2270_ _2648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5652__A1 _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7997_ _0297_ clknet_leaf_37_clk_i memory\[21\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6948_ _1133_ memory\[16\]\[17\] _3444_ _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4758__A3 _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6879_ _3415_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8618_ _0918_ clknet_leaf_88_clk_i memory\[0\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8549_ _0849_ clknet_leaf_117_clk_i memory\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5128__S _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3935__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4032__S _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7343__S _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7180__I1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4967__S _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5891__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5643__A1 _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5597__I _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5946__A2 _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7518__S _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7320__A1 _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3980__I1 _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4230_ _1314_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4161_ _1273_ memory\[15\]\[16\] _1261_ _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6377__B _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6096__C _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5634__A1 _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4092_ _1226_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7920_ _0220_ clknet_leaf_93_clk_i memory\[1\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_132_clk_i_I clknet_4_9_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7851_ _0151_ clknet_leaf_102_clk_i memory\[17\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6802_ _1123_ memory\[9\]\[12\] _3372_ _3375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4994_ memory\[27\]\[13\] _1198_ _1722_ _1726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6985__I1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7782_ _0082_ clknet_leaf_157_clk_i memory\[15\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3945_ net10 _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_15_0_clk_i clknet_0_clk_i clknet_4_15_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_92_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6733_ _1903_ memory\[27\]\[31\] _3318_ _1882_ _3319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_34_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6664_ _1873_ _3251_ _2961_ _3252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5615_ memory\[2\]\[6\] memory\[3\]\[6\] _1992_ _2226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8403_ _0703_ clknet_leaf_32_clk_i memory\[16\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4748__I0 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3876_ _1076_ memory\[7\]\[24\] _1066_ _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6362__A2 _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7227__I _3577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6595_ _2884_ _3184_ _1913_ _3185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8334_ _0634_ clknet_leaf_98_clk_i memory\[9\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5546_ memory\[23\]\[5\] _1896_ _2157_ _1899_ _2158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_131_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4787__S _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_57_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8265_ _0565_ clknet_leaf_126_clk_i memory\[30\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5477_ _1987_ memory\[1\]\[3\] _2090_ _2043_ _2091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3971__I1 _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7216_ _3594_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4428_ _1421_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5173__I0 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7162__I1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8196_ _0496_ clknet_leaf_135_clk_i memory\[28\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7147_ memory\[11\]\[14\] _1200_ _3553_ _3558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4359_ _1384_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_70_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7078_ _3521_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6029_ memory\[16\]\[15\] memory\[17\]\[15\] _2630_ _2631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5625__A1 _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6050__A1 _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7338__S _3650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6041__I _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6105__A2 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7073__S _3517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7153__I1 _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__A1 _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5616__A1 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6644__C _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5919__A2 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7248__S _3577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6344__A2 _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6380_ _1879_ _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5400_ _1871_ _1873_ memory\[25\]\[2\] _2015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5331_ memory\[4\]\[0\] memory\[5\]\[0\] _1935_ _1948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6886__I _3396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8050_ _0350_ clknet_leaf_45_clk_i memory\[23\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4400__S _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5155__I0 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7001_ _3468_ _3480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5262_ _1371_ _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5193_ _1831_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4213_ _1305_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__I0 _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4144_ _1262_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_39_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5231__S _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6280__A1 _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4075_ net19 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_108_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7903_ _0203_ clknet_leaf_182_clk_i memory\[18\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7834_ _0134_ clknet_leaf_12_clk_i memory\[29\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_121_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7765_ _0065_ clknet_leaf_188_clk_i memory\[12\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6716_ _1909_ _3302_ _1994_ _3303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4977_ memory\[27\]\[5\] _1181_ _1711_ _1717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_137_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7696_ _1133_ memory\[7\]\[17\] _1065_ _3848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3928_ _1113_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3859_ _1058_ _1062_ _1064_ _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_62_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6647_ memory\[24\]\[29\] _1858_ _3235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6335__A2 _2930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6997__S _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6578_ _1876_ memory\[19\]\[27\] _3167_ _2003_ _3168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_15_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5529_ _2005_ _2007_ memory\[5\]\[4\] _2142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_42_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8317_ _0617_ clknet_leaf_192_clk_i net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8248_ _0548_ clknet_leaf_204_clk_i memory\[2\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8179_ _0479_ clknet_leaf_44_clk_i memory\[27\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7068__S _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6326__A2 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6700__S _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4220__S _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7126__I1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7531__S _3759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6655__B _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5051__S _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5880_ memory\[30\]\[12\] memory\[31\]\[12\] _2066_ _2485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4890__S _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4900_ _1242_ memory\[26\]\[1\] _1674_ _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6014__A1 _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4831_ _1639_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_134_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7550_ memory\[5\]\[11\] net8 _3770_ _3772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_103_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4762_ memory\[24\]\[0\] _1164_ _1602_ _1603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7481_ _1121_ memory\[10\]\[11\] _3733_ _3735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4693_ _1564_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6501_ memory\[15\]\[25\] _2823_ _3092_ _2773_ _3093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_102_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6432_ _2938_ _2939_ memory\[5\]\[23\] _3026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_125_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6363_ _2674_ memory\[18\]\[22\] _2958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_23_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8102_ _0402_ clknet_leaf_164_clk_i memory\[25\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5128__I0 _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5314_ _1930_ memory\[10\]\[0\] _1931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6294_ _2515_ memory\[7\]\[20\] _2890_ _2517_ _2891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_11_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4130__S _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5828__A1 _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8033_ _0333_ clknet_leaf_165_clk_i memory\[23\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5245_ _1861_ _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5176_ _1822_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4127_ _1250_ memory\[15\]\[5\] _1240_ _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4058_ _1203_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4103__I1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6005__A1 _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6800__I0 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7817_ _0117_ clknet_leaf_127_clk_i memory\[29\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_65_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4305__S _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5628__C _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7748_ _0048_ clknet_leaf_158_clk_i memory\[12\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7679_ _3839_ _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7616__S _3806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5136__S _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7108__I1 _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5119__I0 _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4590__I1 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5819__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4975__S _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7351__S _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6244__A1 _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_179_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5554__B _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3853__I net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6369__C _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5030_ _1744_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6483__A1 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7283__I0 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6981_ memory\[13\]\[0\] _1164_ _3469_ _3470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5932_ memory\[22\]\[13\] _2536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8720_ _1020_ clknet_leaf_70_clk_i memory\[6\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_105_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ memory\[4\]\[11\] _2468_ _2469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8651_ _0951_ clknet_leaf_91_clk_i memory\[10\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5794_ _2163_ _2400_ _2029_ _2401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8582_ _0882_ clknet_leaf_114_clk_i memory\[4\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7602_ _3799_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4814_ memory\[24\]\[25\] _1223_ _1624_ _1630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7533_ memory\[5\]\[3\] net31 _3759_ _3763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4745_ _1591_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_134_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3964__S _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7436__S _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4676_ memory\[22\]\[27\] _1227_ _1546_ _1554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7464_ _1104_ memory\[10\]\[3\] _3722_ _3726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5464__B _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7395_ _3689_ _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6415_ memory\[14\]\[23\] _3009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_116_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4572__I1 _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6346_ _2922_ _2927_ _2932_ _2941_ _2894_ _2942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__4795__S _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8016_ _0316_ clknet_leaf_54_clk_i memory\[22\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6474__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6277_ memory\[15\]\[20\] _2823_ _2873_ _2773_ _2874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5228_ _1849_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input30_I data_i[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5159_ _1154_ memory\[2\]\[27\] _1805_ _1813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_180_clk_i_I clknet_4_9_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7577__I1 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4035__S _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4260__I0 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_209_clk_i clknet_4_2_0_clk_i clknet_leaf_209_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_117_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6701__A2 _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4563__I1 _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7081__S _3517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6768__A2 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7256__S _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ memory\[20\]\[23\] _1219_ _1472_ _1476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4461_ _1074_ memory\[1\]\[23\] _1435_ _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6099__C _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6200_ _1856_ _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7180_ memory\[11\]\[30\] _1233_ _3541_ _3575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6131_ _2313_ _2730_ _2643_ _2731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4392_ _1074_ memory\[18\]\[23\] _1398_ _1402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6062_ _2574_ memory\[28\]\[16\] _2663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6456__B2 _3048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5013_ memory\[27\]\[22\] _1217_ _1733_ _1736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6208__A1 _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7256__I0 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6964_ _3460_ _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5915_ _2467_ _2514_ _2518_ _2519_ _2520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_49_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6895_ memory\[14\]\[24\] _1221_ _3419_ _3424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8703_ _1003_ clknet_leaf_186_clk_i memory\[5\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5846_ memory\[14\]\[11\] _2452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_119_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8634_ _0934_ clknet_leaf_207_clk_i memory\[0\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5777_ _1866_ _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_180_clk_i clknet_4_9_0_clk_i clknet_leaf_180_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_8_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8565_ _0865_ clknet_leaf_201_clk_i memory\[3\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7166__S _3564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8496_ _0796_ clknet_leaf_66_clk_i memory\[11\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4793__I1 _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4728_ _1582_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7516_ _1156_ memory\[10\]\[28\] _3744_ _3753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_127_clk_i_I clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4659_ memory\[22\]\[19\] _1210_ _1535_ _1545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7447_ _3716_ _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6695__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_195_clk_i clknet_4_2_0_clk_i clknet_leaf_195_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_101_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7378_ _1154_ memory\[4\]\[27\] _3672_ _3680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6329_ memory\[8\]\[21\] memory\[9\]\[21\] _2780_ _2925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7495__I0 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5641__C _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6737__C _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_133_clk_i clknet_4_9_0_clk_i clknet_leaf_133_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_94_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5369__B _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_148_clk_i clknet_4_11_0_clk_i clknet_leaf_148_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_137_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4233__I0 _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4536__I1 _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6438__A1 _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5123__I _1782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7238__I0 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3961_ memory\[19\]\[18\] _1135_ _1119_ _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6610__A1 _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5700_ _2305_ _1921_ _2308_ _1927_ _2309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_9_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6680_ _3265_ _3267_ _2887_ _3268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3892_ _1086_ memory\[7\]\[29\] _1087_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5631_ _2108_ memory\[28\]\[7\] _2241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_61_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5562_ _1882_ _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8350_ _0650_ clknet_leaf_169_clk_i memory\[9\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4513_ memory\[20\]\[15\] _1202_ _1461_ _1467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8281_ _0581_ clknet_leaf_17_clk_i memory\[30\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7301_ _3639_ _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7232_ _1144_ memory\[8\]\[22\] _3600_ _3603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6677__A1 _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5493_ _1871_ _2060_ memory\[25\]\[4\] _2106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4444_ _1271_ memory\[1\]\[15\] _1424_ _1430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_113_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4375_ _1271_ memory\[18\]\[15\] _1387_ _1393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7163_ _3566_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6114_ memory\[20\]\[17\] memory\[21\]\[17\] _2346_ _2714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_11_0_clk_i clknet_0_clk_i clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7094_ memory\[31\]\[21\] _1215_ _3528_ _3530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6557__C _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6045_ _2267_ memory\[1\]\[15\] _2646_ _2509_ _2647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5101__A1 _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_50_clk_i clknet_4_5_0_clk_i clknet_leaf_50_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_119_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_53_clk_i_I clknet_4_5_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7996_ _0296_ clknet_leaf_10_clk_i memory\[21\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6601__A1 _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_65_clk_i clknet_4_13_0_clk_i clknet_leaf_65_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_124_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6947_ _3451_ _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4463__I0 _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6878_ memory\[14\]\[16\] _1204_ _3408_ _3415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5829_ _2337_ _2060_ memory\[25\]\[11\] _2435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8617_ _0917_ clknet_leaf_111_clk_i memory\[0\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8548_ _0848_ clknet_leaf_149_clk_i memory\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4766__I1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7624__S _3806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8479_ _0779_ clknet_leaf_180_clk_i memory\[31\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6748__B _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3951__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7468__I0 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6467__C _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output61_I net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4983__S _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_18_clk_i clknet_4_1_0_clk_i clknet_leaf_18_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4782__I _1601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6199__A3 _2795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4206__I0 _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5319__S _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4509__I1 _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6659__B2 _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4160_ net13 _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4091_ memory\[12\]\[26\] _1225_ _1213_ _1226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7850_ _0150_ clknet_leaf_87_clk_i memory\[17\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6801_ _3374_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4993_ _1725_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5398__A1 _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7781_ _0081_ clknet_leaf_157_clk_i memory\[15\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4996__I1 _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3944_ _1124_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6732_ _1935_ memory\[26\]\[31\] _3318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_34_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6663_ memory\[16\]\[29\] memory\[17\]\[29\] _1885_ _3251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3875_ net22 _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8402_ _0702_ clknet_leaf_76_clk_i memory\[16\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5614_ _1987_ memory\[1\]\[6\] _2224_ _2043_ _2225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_14_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4133__S _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5229__S _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6594_ memory\[2\]\[27\] memory\[3\]\[27\] _1911_ _3184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8333_ _0633_ clknet_leaf_98_clk_i memory\[9\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7444__S _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5545_ memory\[20\]\[5\] memory\[21\]\[5\] _1897_ _2157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7698__I0 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8264_ _0564_ clknet_leaf_123_clk_i memory\[30\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5476_ _1988_ memory\[0\]\[3\] _2090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_14_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7215_ _1127_ memory\[8\]\[14\] _3589_ _3594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4427_ _1254_ memory\[1\]\[7\] _1413_ _1421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8195_ _0495_ clknet_leaf_135_clk_i memory\[28\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7146_ _3557_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5873__A2 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4358_ _1254_ memory\[18\]\[7\] _1376_ _1384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_70_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7077_ memory\[31\]\[13\] _1198_ _3517_ _3521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4289_ _1345_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6028_ _1884_ _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5698__I _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4436__I0 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7979_ _0279_ clknet_leaf_49_clk_i memory\[21\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6750__C _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__A1 _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3882__S _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4218__S _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4427__I0 _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7529__S _3759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6660__C _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5049__S _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7264__S _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4888__S _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5330_ _1929_ memory\[7\]\[0\] _1946_ _1932_ _1947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5261_ _1877_ memory\[28\]\[0\] _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_50_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4212_ _1248_ memory\[29\]\[4\] _1300_ _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7000_ _3479_ _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5192_ _1118_ memory\[30\]\[10\] _1830_ _1831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4143_ _1260_ memory\[15\]\[10\] _1261_ _1262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5512__S _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5607__A2 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4074_ _1214_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_39_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7902_ _0202_ clknet_leaf_183_clk_i memory\[18\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_108_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7833_ _0133_ clknet_leaf_12_clk_i memory\[29\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7764_ _0064_ clknet_leaf_27_clk_i memory\[12\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4969__I1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5091__I0 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6715_ memory\[8\]\[30\] memory\[9\]\[30\] _1992_ _3302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4976_ _1716_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5791__A1 _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7695_ _3847_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3927_ memory\[19\]\[7\] _1112_ _1098_ _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3858_ net4 _1063_ _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6646_ _2846_ _3213_ _3233_ _3234_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_116_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6577_ _1877_ memory\[18\]\[27\] _3167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_15_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7174__S _3564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5528_ _2049_ memory\[7\]\[4\] _2140_ _2051_ _2141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_15_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8316_ _0616_ clknet_leaf_18_clk_i net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8247_ _0547_ clknet_leaf_202_clk_i memory\[2\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5459_ _2070_ _1894_ _2072_ _1901_ _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_8178_ _0478_ clknet_leaf_43_clk_i memory\[27\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5930__B _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7129_ _3548_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4038__S _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7349__S _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6023__A2 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7071__I1 _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_175_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6001__B _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7062__I1 _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4830_ _1237_ memory\[25\]\[0\] _1638_ _1639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_44_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_103_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4761_ _1601_ _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_44_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7480_ _3734_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _1242_ memory\[23\]\[1\] _1562_ _1564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6500_ memory\[12\]\[25\] memory\[13\]\[25\] _2919_ _3092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6431_ _2981_ memory\[7\]\[23\] _3024_ _2983_ _3025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_114_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6362_ _2954_ _2760_ _2956_ _2716_ _2957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__5507__S _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5313_ _1869_ _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8101_ _0401_ clknet_leaf_164_clk_i memory\[25\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_54_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5306__I _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6293_ _2562_ memory\[6\]\[20\] _2890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6876__I1 _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8032_ _0332_ clknet_leaf_132_clk_i memory\[22\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5244_ _1295_ _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5175_ _1102_ memory\[30\]\[2\] _1819_ _1822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4126_ net33 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6565__C _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4057_ memory\[12\]\[15\] _1202_ _1192_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6581__B _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6005__A2 _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7816_ _0116_ clknet_leaf_122_clk_i memory\[29\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5064__I0 _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4959_ _1706_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7747_ _0047_ clknet_leaf_159_clk_i memory\[12\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7678_ _1114_ memory\[7\]\[8\] _3837_ _3839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5516__A1 _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6629_ _2828_ memory\[10\]\[28\] _3218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_22_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7632__S _3806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5819__A2 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6492__A2 _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4878__I0 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7431__I _3685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6244__A2 _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7079__S _3517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4007__A1 _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5755__A1 _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5835__B _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4231__S _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4869__I0 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5062__S _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6980_ _3468_ _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5931_ _2531_ _2534_ _2291_ _2535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_105_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4097__I1 _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5994__A1 _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5796__I _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7035__I1 _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8650_ _0950_ clknet_leaf_86_clk_i memory\[10\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4406__S _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5862_ _1858_ _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5793_ memory\[16\]\[10\] memory\[17\]\[10\] _2164_ _2400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8581_ _0881_ clknet_leaf_117_clk_i memory\[4\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7601_ memory\[6\]\[3\] net31 _3795_ _3799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4813_ _1629_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7532_ _3762_ _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4744_ _1080_ memory\[23\]\[26\] _1584_ _1591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6621__S _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5745__B _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4675_ _1553_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7463_ _3725_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6414_ _2993_ _2998_ _3002_ _3007_ _2869_ _3008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_7394_ _1102_ memory\[0\]\[2\] _3686_ _3689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_131_Right_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_116_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3980__S _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6345_ _2933_ _2935_ _2937_ _2940_ _2941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_110_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7452__S _3685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6849__I1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6276_ memory\[12\]\[20\] memory\[13\]\[20\] _2453_ _2873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8015_ _0315_ clknet_leaf_51_clk_i memory\[22\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_47_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5227_ _1154_ memory\[30\]\[27\] _1841_ _1849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6474__A2 _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5480__B _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5158_ _1812_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input23_I data_i[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4109_ _1057_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5089_ _1080_ memory\[28\]\[26\] _1769_ _1776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_123_clk_i_I clknet_4_14_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4088__I1 _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5037__I0 _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4316__S _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_56_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6785__I0 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5655__B _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3954__I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5147__S _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4051__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_48_clk_i_I clknet_4_5_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6217__A2 _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5610__S _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4079__I1 _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5728__A1 _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7537__S _3759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4025__I net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5200__I0 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6153__A1 _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4460_ _1438_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4391_ _1401_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6130_ memory\[8\]\[17\] memory\[9\]\[17\] _2314_ _2730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7272__S _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6061_ _2332_ _2658_ _2660_ _2661_ _2662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_111_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5012_ _1735_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6616__S _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5967__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6963_ _1148_ memory\[16\]\[24\] _3455_ _3460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7008__I1 _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5914_ _2472_ _2473_ memory\[5\]\[12\] _2519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_9_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5459__C _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6894_ _3423_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8702_ _1002_ clknet_leaf_196_clk_i memory\[5\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4136__S _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5719__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5845_ _2436_ _2441_ _2445_ _2450_ _2403_ _2451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_75_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4490__I1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8633_ _0933_ clknet_leaf_207_clk_i memory\[0\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5776_ _1957_ memory\[26\]\[10\] _2383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_90_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8564_ _0864_ clknet_leaf_81_clk_i memory\[3\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5475__B _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8495_ _0795_ clknet_leaf_66_clk_i memory\[11\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4727_ _1277_ memory\[23\]\[18\] _1573_ _1582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7515_ _3752_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6144__A1 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4658_ _1544_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7192__I0 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7446_ _1154_ memory\[0\]\[27\] _3708_ _3716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_130_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4589_ _1507_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7182__S _3541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7377_ _3679_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6328_ _2776_ memory\[11\]\[21\] _2923_ _2640_ _2924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_73_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6259_ _2529_ memory\[29\]\[20\] _2854_ _2855_ _2856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_4_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5430__S _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7357__S _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3885__S _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6383__A1 _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6135__A1 _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_73_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__S _3528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5605__S _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__C _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_82_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3960_ net15 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_86_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3891_ _1065_ _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_72_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5630_ _1857_ _2236_ _2238_ _2239_ _2240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__6374__A1 _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5561_ _1930_ memory\[10\]\[5\] _2173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_5_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4512_ _1466_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_108_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8280_ _0580_ clknet_leaf_3_clk_i memory\[30\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7300_ _1144_ memory\[3\]\[22\] _3636_ _3639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5492_ _1862_ memory\[27\]\[4\] _2104_ _1867_ _2105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6126__B2 _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7231_ _3602_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4443_ _1429_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_113_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6921__I0 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4374_ _1392_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7162_ memory\[11\]\[21\] _1215_ _3564_ _3566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6113_ _1061_ _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7093_ _3529_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6429__A2 _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6044_ _2318_ memory\[0\]\[15\] _2646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_119_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_208_clk_i clknet_4_2_0_clk_i clknet_leaf_208_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7995_ _0295_ clknet_leaf_40_clk_i memory\[21\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6946_ _1131_ memory\[16\]\[16\] _3444_ _3451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_124_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6877_ _3414_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6081__S _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5828_ _2382_ memory\[27\]\[11\] _2433_ _2384_ _2434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_107_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8616_ _0916_ clknet_leaf_112_clk_i memory\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5759_ _2364_ _2366_ _1939_ _2367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8547_ _0847_ clknet_leaf_152_clk_i memory\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8478_ _0778_ clknet_leaf_20_clk_i memory\[31\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7429_ _1137_ memory\[0\]\[19\] _3697_ _3707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_9_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5340__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6764__B _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output54_I net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7087__S _3517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6108__A1 _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5843__B _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6659__A2 _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7320__A3 _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4390__I0 _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7550__S _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6674__B _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4090_ net24 _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5070__S _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6800_ _1121_ memory\[9\]\[11\] _3372_ _3374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4992_ memory\[27\]\[12\] _1196_ _1722_ _1725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_81_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6595__A1 _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_194_clk_i clknet_4_2_0_clk_i clknet_leaf_194_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7780_ _0080_ clknet_leaf_157_clk_i memory\[15\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3943_ memory\[19\]\[12\] _1123_ _1119_ _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_105_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6731_ memory\[24\]\[31\] _1858_ _3317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_34_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6662_ _1876_ memory\[19\]\[29\] _3249_ _2003_ _3250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_46_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3874_ _1075_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6347__A1 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8401_ _0701_ clknet_leaf_70_clk_i memory\[16\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5613_ _1988_ memory\[0\]\[6\] _2224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_61_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8332_ _0632_ clknet_leaf_97_clk_i memory\[9\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6593_ _1904_ memory\[1\]\[27\] _3182_ _2975_ _3183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_5_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5544_ memory\[22\]\[5\] _2156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_124_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8263_ _0563_ clknet_leaf_123_clk_i memory\[30\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_132_clk_i clknet_4_9_0_clk_i clknet_leaf_132_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5475_ _2086_ _2088_ _1939_ _2089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7214_ _3593_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4426_ _1420_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8194_ _0494_ clknet_leaf_130_clk_i memory\[28\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5472__C _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7145_ memory\[11\]\[13\] _1198_ _3553_ _3557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4381__I0 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4357_ _1383_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_70_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7460__S _3722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7076_ _3520_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4288_ _1256_ memory\[17\]\[8\] _1336_ _1345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_147_clk_i clknet_4_11_0_clk_i clknet_leaf_147_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6076__S _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6027_ _1872_ _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4133__I0 _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4684__I1 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_9_0_clk_i clknet_0_clk_i clknet_4_9_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6804__S _3372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7622__I1 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7978_ _0278_ clknet_leaf_131_clk_i memory\[21\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6929_ _1114_ memory\[16\]\[8\] _3433_ _3442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5647__C _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4324__S _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7386__I0 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6759__B _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5663__B _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5155__S _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4994__S _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7370__S _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7310__I0 _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4124__I0 _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_171_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7613__I1 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6577__A1 _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7545__S _3759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3872__I net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5260_ _1863_ _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_51_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_64_clk_i clknet_4_7_0_clk_i clknet_leaf_64_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_96_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4211_ _1304_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6501__B2 _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5191_ _1818_ _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_10_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5799__I _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4142_ _1239_ _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4115__I0 _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4073_ memory\[12\]\[20\] _1212_ _1213_ _1214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_39_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_79_clk_i clknet_4_6_0_clk_i clknet_leaf_79_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4666__I1 _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7901_ _0201_ clknet_leaf_184_clk_i memory\[18\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_108_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7832_ _0132_ clknet_leaf_13_clk_i memory\[29\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6568__A1 _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7763_ _0063_ clknet_leaf_75_clk_i memory\[12\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4975_ memory\[27\]\[4\] _1179_ _1711_ _1716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3926_ net35 _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_86_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6714_ _1987_ memory\[11\]\[30\] _3300_ _1907_ _3301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_128_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7694_ _1131_ memory\[7\]\[16\] _3837_ _3847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7368__I0 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_clk_i clknet_4_1_0_clk_i clknet_leaf_17_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3983__S _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6645_ _1854_ net59 _3234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3857_ net5 _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_117_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6576_ _3163_ _2760_ _3165_ _1937_ _3166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_61_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5527_ _2096_ memory\[6\]\[4\] _2140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8315_ _0615_ clknet_leaf_17_clk_i net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8246_ _0546_ clknet_leaf_202_clk_i memory\[2\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6298__C _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4354__I0 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5458_ memory\[23\]\[3\] _1896_ _2071_ _1899_ _2072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8177_ _0477_ clknet_leaf_48_clk_i memory\[27\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5389_ _1870_ _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7190__S _3578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4409_ _1410_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7128_ memory\[11\]\[5\] _1181_ _3542_ _3548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7059_ _3511_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4657__I1 _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A1 _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6761__C _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4054__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3957__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7359__I0 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5534__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_118_clk_i_I clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4229__S _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4028__I net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6444__S _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_103_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _1600_ _1601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4820__I1 _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7275__S _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4691_ _1563_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _1864_ memory\[6\]\[23\] _3024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_125_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6361_ memory\[23\]\[22\] _2713_ _2955_ _2671_ _2956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_24_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5312_ _1903_ _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8100_ _0400_ clknet_leaf_176_clk_i memory\[25\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5289__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6292_ memory\[4\]\[20\] _2468_ _2889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7522__I0 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8031_ _0331_ clknet_leaf_132_clk_i memory\[22\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4336__I0 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5243_ memory\[24\]\[0\] _1859_ _1860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5174_ _1821_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4125_ _1249_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4139__S _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5322__I _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4056_ net12 _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_79_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7815_ _0115_ clknet_leaf_128_clk_i memory\[29\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_65_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4958_ _1086_ memory\[26\]\[29\] _1696_ _1706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7746_ _0046_ clknet_leaf_156_clk_i memory\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7677_ _3838_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4889_ _1669_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3909_ memory\[19\]\[1\] _1100_ _1098_ _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6713__A1 _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6628_ _3214_ _2872_ _3216_ _2826_ _3217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_117_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6559_ _2933_ _3146_ _3148_ _3149_ _3150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__5941__B _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8229_ _0529_ clknet_leaf_117_clk_i memory\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6756__C _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3888__S _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6264__S _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_44_clk_i_I clknet_4_4_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4007__A2 _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7159__I _3541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6704__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7504__I0 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4318__I0 _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6666__C _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_49_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5930_ _2288_ _2533_ _2200_ _2534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_105_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7600_ _3798_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ _1058_ _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5792_ _2160_ memory\[19\]\[10\] _2398_ _2075_ _2399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8580_ _0880_ clknet_leaf_118_clk_i memory\[4\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4812_ memory\[24\]\[24\] _1221_ _1624_ _1629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7531_ memory\[5\]\[2\] net28 _3759_ _3762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4743_ _1590_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7462_ _1102_ memory\[10\]\[2\] _3722_ _3725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4674_ memory\[22\]\[26\] _1225_ _1546_ _1553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6413_ _3004_ _3006_ _2768_ _3007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_113_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5317__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7393_ _3688_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6344_ _2938_ _2939_ memory\[5\]\[21\] _2940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_101_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4309__I0 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6275_ _1893_ _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8014_ _0314_ clknet_leaf_54_clk_i memory\[22\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_102_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6576__C _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5226_ _1848_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5157_ _1152_ memory\[2\]\[26\] _1805_ _1812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4108_ net6 _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5088_ _1775_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input16_I data_i[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4039_ _1190_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6812__S _3372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7729_ _0029_ clknet_leaf_72_clk_i memory\[19\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4332__S _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7643__S _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5163__S _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3970__I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5673__A1 _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4507__S _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5425__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4041__I _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ _1072_ memory\[18\]\[22\] _1398_ _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_0_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input8_I data_i[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6060_ _2337_ _2526_ memory\[25\]\[16\] _2661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_111_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4711__I0 _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5011_ memory\[27\]\[21\] _1215_ _1733_ _1735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4417__S _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6962_ _3459_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5913_ _2515_ memory\[7\]\[12\] _2516_ _2517_ _2518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_75_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6893_ memory\[14\]\[23\] _1219_ _3419_ _3423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8701_ _1001_ clknet_leaf_194_clk_i memory\[5\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5019__I1 _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5844_ _2447_ _2449_ _2302_ _2450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_62_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8632_ _0932_ clknet_leaf_193_clk_i memory\[0\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8563_ _0863_ clknet_leaf_83_clk_i memory\[3\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4152__S _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5775_ _1861_ _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7514_ _1154_ memory\[10\]\[27\] _3744_ _3752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8494_ _0794_ clknet_leaf_94_clk_i memory\[11\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4726_ _1581_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4657_ memory\[22\]\[18\] _1208_ _1535_ _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7445_ _3715_ _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7376_ _1152_ memory\[4\]\[26\] _3672_ _3679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4588_ memory\[21\]\[18\] _1208_ _1498_ _1507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3902__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6327_ _2828_ memory\[10\]\[21\] _2923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4950__I0 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5655__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6258_ _1879_ _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5209_ _1839_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6189_ _2418_ _2787_ _2602_ _2788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4702__I0 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_217_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4126__I net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6542__S _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3992__I1 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5194__I0 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6497__B _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4237__S _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6997__I1 _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__B2 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7548__S _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3890_ net27 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5068__S _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3875__I net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5560_ _2169_ _1921_ _2171_ _1927_ _2172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4511_ memory\[20\]\[14\] _1200_ _1461_ _1466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_102_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6126__A2 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3983__I1 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5491_ _1957_ memory\[26\]\[4\] _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7283__S _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4442_ _1269_ memory\[1\]\[14\] _1424_ _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5185__I0 _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7230_ _1142_ memory\[8\]\[21\] _3600_ _3602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4700__S _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7174__I1 _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_166_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5885__B2 _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4373_ _1269_ memory\[18\]\[14\] _1387_ _1392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7161_ _3565_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6112_ memory\[22\]\[17\] _2712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7092_ memory\[31\]\[20\] _1212_ _3528_ _3529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6043_ _2641_ _2644_ _2414_ _2645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_1_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7994_ _0294_ clknet_leaf_40_clk_i memory\[21\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6945_ _3450_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6062__A1 _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__S _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7458__S _3722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6876_ memory\[14\]\[15\] _1202_ _3408_ _3414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5827_ _2432_ memory\[26\]\[11\] _2433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8615_ _0915_ clknet_leaf_112_clk_i memory\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5758_ _2313_ _2365_ _2177_ _2366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6161__I _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8546_ _0846_ clknet_leaf_152_clk_i memory\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6117__A2 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4709_ _1572_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3974__I1 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8477_ _0777_ clknet_leaf_191_clk_i memory\[31\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5706__S _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5689_ _2208_ memory\[18\]\[8\] _2298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7428_ _3706_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_75_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5876__A1 _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_5_0_clk_i clknet_0_clk_i clknet_4_5_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_102_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4923__I0 _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6110__B _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7359_ _1135_ memory\[4\]\[18\] _3661_ _3670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6537__S _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5628__A1 _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output47_I net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4057__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5240__I _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6053__A1 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7368__S _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6004__C _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5167__I0 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6903__I1 _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4914__I0 _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5619__A1 _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6044__A1 _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_92_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4991_ _1724_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6182__S _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _1954_ _3295_ _3315_ _3316_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3942_ net9 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_34_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6661_ _1877_ memory\[18\]\[29\] _3249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6347__A2 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3873_ _1074_ memory\[7\]\[23\] _1066_ _1075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8400_ _0700_ clknet_leaf_70_clk_i memory\[16\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5612_ _2220_ _2222_ _1939_ _2223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_14_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6592_ _2784_ memory\[0\]\[27\] _3182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8331_ _0631_ clknet_leaf_90_clk_i memory\[9\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5543_ _2152_ _2154_ _1890_ _2155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7147__I1 _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8262_ _0562_ clknet_leaf_122_clk_i memory\[30\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5474_ _1934_ _2087_ _1937_ _2088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5753__C _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7213_ _1125_ memory\[8\]\[13\] _3589_ _3593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4425_ _1252_ memory\[1\]\[6\] _1413_ _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8193_ _0493_ clknet_leaf_135_clk_i memory\[28\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7144_ _3556_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4356_ _1252_ memory\[18\]\[6\] _1376_ _1383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7075_ memory\[31\]\[12\] _1196_ _3517_ _3520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4287_ _1344_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6026_ _2626_ memory\[19\]\[15\] _2627_ _2541_ _2628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6035__B2 _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3892__I0 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7977_ _0277_ clknet_leaf_129_clk_i memory\[21\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7188__S _3578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6586__A2 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6928_ _3441_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__S _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6859_ memory\[14\]\[7\] _1185_ _3397_ _3405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8529_ _0829_ clknet_leaf_97_clk_i memory\[8\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5149__I0 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5849__B2 _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7651__S _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5171__S _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6494__C _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_114_clk_i_I clknet_4_15_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6026__A1 _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7098__S _3528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6821__I0 _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4515__S _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_99_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5854__B _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_207_clk_i clknet_4_2_0_clk_i clknet_leaf_207_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4250__S _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_clk_i_I clknet_4_4_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4210_ _1246_ memory\[29\]\[3\] _1300_ _1304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6501__A2 _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _1829_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4141_ net7 _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_0_clk_i clk_i clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5081__S _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6265__B2 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4072_ _1170_ _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_39_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7900_ _0200_ clknet_leaf_184_clk_i memory\[18\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6905__S _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6812__I0 _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7831_ _0131_ clknet_leaf_22_clk_i memory\[29\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4425__S _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7762_ _0062_ clknet_leaf_75_clk_i memory\[12\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4974_ _1715_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7693_ _3846_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3925_ _1111_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6713_ _1988_ memory\[10\]\[30\] _3300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_129_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4224__I _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6644_ _3217_ _3222_ _3227_ _3232_ _2894_ _3233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_117_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5764__B _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3856_ net38 _1061_ _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_62_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6575_ memory\[23\]\[27\] _1895_ _3164_ _2006_ _3165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5526_ memory\[4\]\[4\] _1998_ _2139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8314_ _0614_ clknet_leaf_17_clk_i net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8245_ _0545_ clknet_leaf_201_clk_i memory\[2\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5457_ memory\[20\]\[3\] memory\[21\]\[3\] _1897_ _2071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5055__I _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4408_ _1091_ memory\[18\]\[31\] _1375_ _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8176_ _0476_ clknet_leaf_48_clk_i memory\[27\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5388_ _2000_ memory\[7\]\[1\] _2002_ _2003_ _2004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6595__B _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4339_ _1059_ _1371_ _1372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7127_ _3547_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7058_ memory\[31\]\[4\] _1179_ _3506_ _3511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6256__A1 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4106__I1 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6009_ _2380_ _2589_ _2610_ _2611_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_97_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6008__A1 _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4290__I0 _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6731__A2 _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3973__I net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4593__I1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_40_clk_i_I clknet_4_4_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_193_clk_i clknet_4_2_0_clk_i clknet_leaf_193_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_130_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6247__A1 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5470__A2 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_131_clk_i clknet_4_12_0_clk_i clknet_leaf_131_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_16_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7556__S _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4044__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_146_clk_i clknet_4_11_0_clk_i clknet_leaf_146_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4690_ _1237_ memory\[23\]\[0\] _1562_ _1563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4584__I1 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6360_ memory\[20\]\[22\] memory\[21\]\[22\] _2812_ _2955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5311_ _1920_ _1921_ _1926_ _1927_ _1928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_122_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7291__S _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8030_ _0330_ clknet_leaf_30_clk_i memory\[22\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6291_ _2883_ _2886_ _2887_ _2888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_54_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5242_ _1858_ _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5173_ _1100_ memory\[30\]\[1\] _1819_ _1821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4124_ _1248_ memory\[15\]\[4\] _1240_ _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput1 address_i[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4055_ _1201_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__B _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4155__S _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7814_ _0114_ clknet_leaf_122_clk_i memory\[29\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7589__I1 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6410__A1 _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4272__I0 _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4957_ _1705_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7745_ _0045_ clknet_leaf_150_clk_i memory\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7466__S _3722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7676_ _1112_ memory\[7\]\[7\] _3837_ _3838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3908_ net17 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_62_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4888_ _1084_ memory\[25\]\[28\] _1660_ _1669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6627_ memory\[15\]\[28\] _2823_ _3215_ _1899_ _3216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_105_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6558_ _2938_ _2939_ memory\[5\]\[26\] _3149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_120_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6489_ memory\[22\]\[25\] _3081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5509_ _2119_ _2121_ _1916_ _2122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6477__A1 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8228_ _0528_ clknet_leaf_149_clk_i memory\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8159_ _0459_ clknet_leaf_183_clk_i memory\[26\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7277__I0 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4129__I net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5388__C _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6401__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_63_clk_i clknet_4_7_0_clk_i clknet_leaf_63_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7376__S _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_78_clk_i clknet_4_6_0_clk_i clknet_leaf_78_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6012__C _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7268__I0 _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_16_clk_i clknet_4_1_0_clk_i clknet_leaf_16_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_49_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5443__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6640__A1 _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5860_ _2463_ _2465_ _2421_ _2466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_105_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3878__I net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4811_ _1628_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7440__I0 _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5791_ _2208_ memory\[18\]\[10\] _2398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4254__I0 _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4742_ _1078_ memory\[23\]\[25\] _1584_ _1590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7530_ _3761_ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4673_ _1552_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7461_ _3724_ _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4502__I _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6412_ _2629_ _3005_ _2961_ _3006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7392_ _1100_ memory\[0\]\[1\] _3686_ _3688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4557__I1 _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6343_ _2006_ _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_110_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5761__C _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6459__B2 _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6274_ memory\[14\]\[20\] _2871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8013_ _0313_ clknet_leaf_53_clk_i memory\[22\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5225_ _1152_ memory\[30\]\[26\] _1841_ _1848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5333__I _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3989__S _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5156_ _1811_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5087_ _1078_ memory\[28\]\[25\] _1769_ _1775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6365__S _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4107_ _1236_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4038_ memory\[12\]\[9\] _1189_ _1171_ _1190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_8_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5989_ memory\[15\]\[14\] _2357_ _2591_ _2307_ _2592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__7196__S _3578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7728_ _0028_ clknet_leaf_71_clk_i memory\[19\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4613__S _1486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4412__I _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7659_ memory\[6\]\[31\] net30 _3794_ _3829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_213_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6767__C _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6622__A1 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6007__C _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4787__I1 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7489__I0 _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6677__C _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6249__I _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5010_ _1734_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5664__A2 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_4_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7661__I0 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6613__A1 _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6961_ _1146_ memory\[16\]\[23\] _3455_ _3459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_162_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__I0 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8700_ _1000_ clknet_leaf_3_clk_i memory\[5\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5912_ _1866_ _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6913__S _3433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6892_ _3422_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7413__I0 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5843_ _2163_ _2448_ _2029_ _2449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4227__I0 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8631_ _0931_ clknet_leaf_203_clk_i memory\[0\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5756__C _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8562_ _0862_ clknet_leaf_84_clk_i memory\[3\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_62_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4778__I1 _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5774_ memory\[24\]\[10\] _2333_ _2381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7513_ _3751_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8493_ _0793_ clknet_leaf_94_clk_i memory\[11\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4725_ _1275_ memory\[23\]\[17\] _1573_ _1581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4656_ _1543_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7444_ _1152_ memory\[0\]\[26\] _3708_ _3715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4587_ _1506_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7375_ _3678_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3902__A2 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6326_ _2918_ _2872_ _2921_ _2826_ _2922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_clkbuf_leaf_87_clk_i_I clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6257_ _2574_ memory\[28\]\[20\] _2854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6188_ memory\[2\]\[18\] memory\[3\]\[18\] _2736_ _2787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5208_ _1135_ memory\[30\]\[18\] _1830_ _1839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5139_ _1802_ _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_1_0_clk_i clknet_0_clk_i clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_95_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6823__S _3383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7404__I0 _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4218__I0 _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5666__C _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__I _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4142__I _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6540__B1 _3125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5343__A1 _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5701__I _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_121_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6018__B _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4457__I0 _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__A2 _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7564__S _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5582__A1 _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_130_Left_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4510_ _1465_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_124_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5490_ memory\[24\]\[4\] _1859_ _2103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4441_ _1428_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_109_clk_i_I clknet_4_15_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3891__I _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4987__I _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5885__A2 _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7160_ memory\[11\]\[20\] _1212_ _3564_ _3565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7363__I _3649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4372_ _1391_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6111_ _2708_ _2710_ _2291_ _2711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_59_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5812__S _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7091_ _3505_ _3528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_10_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6042_ _2313_ _2642_ _2643_ _2644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4696__I0 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4448__I0 _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7993_ _0293_ clknet_leaf_40_clk_i memory\[21\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6944_ _1129_ memory\[16\]\[15\] _3444_ _3450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6875_ _3413_ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8614_ _0914_ clknet_leaf_113_clk_i memory\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5826_ _1910_ _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_9_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5757_ memory\[8\]\[9\] memory\[9\]\[9\] _2314_ _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7474__S _3722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8545_ _0845_ clknet_leaf_139_clk_i memory\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4708_ _1258_ memory\[23\]\[9\] _1562_ _1572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8476_ _0776_ clknet_leaf_4_clk_i memory\[31\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7427_ _1135_ memory\[0\]\[18\] _3697_ _3706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5688_ _2293_ _2294_ _2296_ _2250_ _2297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_75_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5325__A1 _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4897__I _1673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5876__A2 _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4639_ _1534_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_9_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7358_ _3669_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7289_ _1133_ memory\[3\]\[17\] _3625_ _3633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6309_ memory\[30\]\[21\] memory\[31\]\[21\] _2532_ _2905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_86_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7649__S _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3976__I net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4073__S _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7384__S _3649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4801__S _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_110_clk_i_I clknet_4_15_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5316__A1 _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_128_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6292__A2 _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4248__S _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4047__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__I1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6463__S _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4990_ memory\[27\]\[11\] _1194_ _1722_ _1724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_35_clk_i_I clknet_4_4_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3941_ _1122_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5079__S _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6660_ _3245_ _1893_ _3247_ _1937_ _3248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3872_ net21 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_128_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5611_ _1934_ _2221_ _2177_ _2222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6591_ _3178_ _3180_ _2880_ _3181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4711__S _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8330_ _0630_ clknet_leaf_89_clk_i memory\[9\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5542_ _1883_ _2153_ _1887_ _2154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6211__B _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ memory\[8\]\[3\] memory\[9\]\[3\] _1935_ _2087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8261_ _0561_ clknet_leaf_120_clk_i memory\[30\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7212_ _3592_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4424_ _1419_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8192_ _0492_ clknet_leaf_134_clk_i memory\[27\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7143_ memory\[11\]\[12\] _1196_ _3553_ _3556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4355_ _1382_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7074_ _3519_ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_70_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4286_ _1254_ memory\[17\]\[7\] _1336_ _1344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4158__S _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6025_ _2208_ memory\[18\]\[15\] _2627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5341__I _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6035__A2 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7083__I1 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7976_ _0276_ clknet_leaf_140_clk_i memory\[21\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5794__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6927_ _1112_ memory\[16\]\[7\] _3433_ _3441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6858_ _3404_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5809_ _2318_ memory\[0\]\[10\] _2416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_107_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6743__B1 _3328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5546__B2 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8528_ _0828_ clknet_leaf_96_clk_i memory\[8\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6789_ _1110_ memory\[9\]\[6\] _3361_ _3368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6121__B _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8459_ _0759_ clknet_leaf_73_clk_i memory\[31\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5849__A2 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6897__I1 _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5085__I0 _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5785__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4832__I0 _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4060__I1 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__B _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6458__S _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4140_ _1259_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6265__A2 _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ net18 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7289__S _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4706__S _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7830_ _0130_ clknet_leaf_14_clk_i memory\[29\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7761_ _0061_ clknet_leaf_58_clk_i memory\[12\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5776__A1 _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4973_ memory\[27\]\[3\] _1177_ _1711_ _1715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7692_ _1129_ memory\[7\]\[15\] _3837_ _3846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3924_ memory\[19\]\[6\] _1110_ _1098_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6921__S _3433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6712_ _3296_ _1894_ _3298_ _1901_ _3299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_129_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5528__A1 _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6643_ _2933_ _3228_ _3230_ _3231_ _3232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_117_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3855_ _1059_ _1060_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4051__I1 _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6574_ memory\[20\]\[27\] memory\[21\]\[27\] _2812_ _3164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4200__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5525_ _2134_ _2137_ _1950_ _2138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_70_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8313_ _0613_ clknet_leaf_18_clk_i net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_119_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8244_ _0544_ clknet_leaf_82_clk_i memory\[2\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5456_ memory\[22\]\[3\] _2070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_100_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4407_ _1409_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8175_ _0475_ clknet_leaf_50_clk_i memory\[27\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5387_ _1866_ _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4338_ _1060_ _1371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_7126_ memory\[11\]\[4\] _1179_ _3542_ _3547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7057_ _3510_ _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4269_ _1334_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6008_ _2330_ net44 _2611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7056__I1 _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A1 _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7959_ _0259_ clknet_leaf_41_clk_i memory\[20\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__S _3383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5955__B _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4042__I1 _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6192__A1 _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5674__C _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5246__I _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6247__A2 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_208_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5058__I0 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4526__S _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5758__A1 _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5357__S _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7636__I _3794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6183__A1 _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5930__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6290_ _1915_ _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5310_ _1058_ _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__6188__S _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5241_ _1168_ _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_54_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5172_ _1820_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4123_ net32 _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4054_ memory\[12\]\[14\] _1200_ _1192_ _1201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput2 address_i[1] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5997__A1 _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4436__S _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5049__I0 _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7813_ _0113_ clknet_leaf_129_clk_i memory\[29\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7744_ _0044_ clknet_leaf_181_clk_i memory\[19\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _1084_ memory\[26\]\[28\] _1696_ _1705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7675_ _1065_ _3837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4887_ _1668_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3907_ _1099_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5221__I0 _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6626_ memory\[12\]\[28\] memory\[13\]\[28\] _2919_ _3215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5921__A1 _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6557_ _2981_ memory\[7\]\[26\] _3147_ _2983_ _3148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5508_ _1909_ _2120_ _2029_ _2121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_4_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6488_ _3077_ _3079_ _2757_ _3080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_157_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5439_ _1997_ _2048_ _2052_ _2053_ _2054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_8227_ _0527_ clknet_leaf_151_clk_i memory\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6477__A2 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8158_ _0458_ clknet_leaf_15_clk_i memory\[26\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6229__A2 _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7109_ _3537_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8089_ _0389_ clknet_leaf_9_clk_i memory\[24\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5669__C _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_206_clk_i clknet_4_2_0_clk_i clknet_leaf_206_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7029__I1 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4346__S _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4145__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7657__S _3794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5177__S _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6165__A1 _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7392__S _3686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5704__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4479__A1 _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5979__B2 _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4256__S _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__I0 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4810_ memory\[24\]\[23\] _1219_ _1624_ _1628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_29_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5790_ _2394_ _2294_ _2396_ _2250_ _2397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_68_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4741_ _1589_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5087__S _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3894__I net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4672_ memory\[22\]\[25\] _1223_ _1546_ _1552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7460_ _1100_ memory\[10\]\[1\] _3722_ _3724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5903__A1 _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6411_ memory\[16\]\[23\] memory\[17\]\[23\] _2630_ _3005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_102_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7391_ _3687_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_116_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6342_ _1870_ _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_110_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6273_ _2853_ _2859_ _2863_ _2868_ _2869_ _2870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_11_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6459__A2 _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8012_ _0312_ clknet_leaf_54_clk_i memory\[22\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5224_ _1847_ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4190__I0 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5155_ _1150_ memory\[2\]\[25\] _1805_ _1811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5086_ _1774_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_16_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4106_ memory\[12\]\[31\] _1235_ _1170_ _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4037_ net37 _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_67_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_83_clk_i_I clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5988_ memory\[12\]\[14\] memory\[13\]\[14\] _2453_ _2591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_192_clk_i clknet_4_3_0_clk_i clknet_leaf_192_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7727_ _0027_ clknet_leaf_89_clk_i memory\[19\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4939_ _1673_ _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6147__A1 _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6180__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7658_ _3828_ _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_133_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6609_ _2798_ _3194_ _3196_ _3197_ _3198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6942__I0 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7589_ memory\[5\]\[30\] net29 _3758_ _3792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_130_clk_i clknet_4_12_0_clk_i clknet_leaf_130_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_7_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_145_clk_i clknet_4_11_0_clk_i clknet_leaf_145_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3979__I net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5399__C _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4076__S _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4484__I1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4804__S _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_43_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6138__A1 _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_11_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6023__C _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6689__A2 _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7186__I0 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5434__I _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6310__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4172__I0 _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6960_ _3458_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_105_clk_i_I clknet_4_15_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5911_ _2096_ memory\[6\]\[12\] _2516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_4_8_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6891_ memory\[14\]\[22\] _1217_ _3419_ _3422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5842_ memory\[16\]\[11\] memory\[17\]\[11\] _2164_ _2448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6377__A1 _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8630_ _0930_ clknet_leaf_194_clk_i memory\[0\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8561_ _0861_ clknet_leaf_93_clk_i memory\[3\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5773_ _1854_ _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_75_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6129__A1 _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4724_ _1580_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7512_ _1152_ memory\[10\]\[26\] _3744_ _3751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8492_ _0792_ clknet_leaf_93_clk_i memory\[11\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4655_ memory\[22\]\[17\] _1206_ _1535_ _1543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5545__S _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7443_ _3714_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4586_ memory\[21\]\[17\] _1206_ _1498_ _1506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7374_ _1150_ memory\[4\]\[25\] _3672_ _3678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6325_ memory\[15\]\[21\] _2823_ _2920_ _2773_ _2921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3902__A3 _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_62_clk_i clknet_4_7_0_clk_i clknet_leaf_62_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6256_ _2798_ _2847_ _2851_ _2852_ _2853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5207_ _1838_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6187_ _2733_ memory\[1\]\[18\] _2785_ _2509_ _2786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6376__S _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5138_ _1275_ memory\[2\]\[17\] _1794_ _1802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_4_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input21_I data_i[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6108__C _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5069_ _1765_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_77_clk_i clknet_4_12_0_clk_i clknet_leaf_77_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_88_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4624__S _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6915__I0 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_clk_i clknet_4_1_0_clk_i clknet_leaf_15_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_105_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6540__B2 _3130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5254__I _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7340__I0 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7643__I1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5857__C _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4534__S _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4440_ _1267_ memory\[1\]\[13\] _1424_ _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_31_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4371_ _1267_ memory\[18\]\[13\] _1387_ _1391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6110_ _2288_ _2709_ _2666_ _2710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_59_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7090_ _3527_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6041_ _1238_ _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_1_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7634__I1 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7992_ _0292_ clknet_leaf_41_clk_i memory\[21\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6598__A1 _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6943_ _3449_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4444__S _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6874_ memory\[14\]\[14\] _1200_ _3408_ _3413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5767__C _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7398__I0 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5825_ memory\[24\]\[11\] _2333_ _2431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8613_ _0913_ clknet_leaf_123_clk_i memory\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5573__A2 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5756_ _2310_ memory\[11\]\[9\] _2363_ _2174_ _2364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_45_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8544_ _0844_ clknet_leaf_168_clk_i memory\[8\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4620__I1 _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5687_ memory\[23\]\[8\] _2247_ _2295_ _2205_ _2296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4707_ _1571_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8475_ _0775_ clknet_leaf_3_clk_i memory\[31\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7426_ _3705_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4638_ memory\[22\]\[9\] _1189_ _1524_ _1534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_75_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6522__A1 _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7357_ _1133_ memory\[4\]\[17\] _3661_ _3669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4569_ memory\[21\]\[9\] _1189_ _1487_ _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7288_ _3632_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7322__I0 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6308_ _2529_ memory\[29\]\[21\] _2903_ _2855_ _2904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6239_ _2418_ _2836_ _2602_ _2837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4136__I0 _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4354__S _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5261__A1 _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7665__S _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5249__I _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6761__A1 _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4611__I1 _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5185__S _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4375__I0 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4127__I0 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4678__I1 _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7616__I1 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3940_ memory\[19\]\[11\] _1121_ _1119_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5587__C _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4264__S _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7575__S _3781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3871_ _1073_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5610_ memory\[8\]\[6\] memory\[9\]\[6\] _1935_ _2221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6590_ _2779_ _3179_ _1994_ _3180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5541_ memory\[30\]\[5\] memory\[31\]\[5\] _2066_ _2153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_14_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8260_ _0560_ clknet_leaf_121_clk_i memory\[30\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5095__S _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7211_ _1123_ memory\[8\]\[12\] _3589_ _3592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5472_ _1929_ memory\[11\]\[3\] _2085_ _1932_ _2086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6504__A1 _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4423_ _1250_ memory\[1\]\[5\] _1413_ _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8191_ _0491_ clknet_leaf_183_clk_i memory\[27\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6919__S _3433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7142_ _3555_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4354_ _1250_ memory\[18\]\[5\] _1376_ _1382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7304__I0 _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7073_ memory\[31\]\[11\] _1194_ _3517_ _3519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_70_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4118__I0 _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4285_ _1343_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6024_ _1861_ _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5491__A1 _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7607__I1 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6654__S _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7975_ _0275_ clknet_leaf_155_clk_i memory\[21\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6926_ _3440_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5497__C _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4174__S _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7485__S _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ memory\[14\]\[6\] _1183_ _3397_ _3404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5808_ _2411_ _2413_ _2414_ _2415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6788_ _3367_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5546__A2 _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4902__S _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8527_ _0827_ clknet_leaf_98_clk_i memory\[8\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5739_ memory\[20\]\[9\] memory\[21\]\[9\] _2346_ _2347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6743__B2 _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8458_ _0758_ clknet_leaf_82_clk_i memory\[31\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7409_ _3696_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8389_ _0689_ clknet_leaf_144_clk_i memory\[16\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6829__S _3383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5960__C _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output52_I net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4148__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6734__A1 _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5537__A2 _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4812__S _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_204_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6498__B1 _3084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4348__I0 _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5870__C _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4070_ _1211_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_39_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_108_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3897__I net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7760_ _0060_ clknet_leaf_61_clk_i memory\[12\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_121_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4972_ _1714_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_121_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3923_ net34 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7691_ _3845_ _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6711_ memory\[15\]\[30\] _1896_ _3297_ _1899_ _3298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_117_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3854_ net2 _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6642_ _2938_ _2939_ memory\[5\]\[28\] _3231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6725__A1 _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6222__B _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6573_ memory\[22\]\[27\] _3163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8312_ _0612_ clknet_leaf_18_clk_i net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5524_ _1941_ _2135_ _2136_ _2137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8243_ _0543_ clknet_leaf_82_clk_i memory\[2\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5455_ _2065_ _2068_ _1890_ _2069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8174_ _0474_ clknet_leaf_47_clk_i memory\[27\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5000__I1 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5553__S _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4406_ _1089_ memory\[18\]\[30\] _1375_ _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7125_ _3546_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5386_ _2001_ memory\[6\]\[1\] _2002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5700__A2 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4169__S _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4337_ _1370_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7056_ memory\[31\]\[3\] _1177_ _3506_ _3510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4268_ _1091_ memory\[29\]\[31\] _1299_ _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6007_ _2593_ _2598_ _2604_ _2609_ _2428_ _2610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__5464__A1 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4199_ _1295_ _1060_ _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_0_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_153_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7958_ _0258_ clknet_leaf_42_clk_i memory\[20\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7889_ _0189_ clknet_leaf_72_clk_i memory\[18\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4814__I1 _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6909_ memory\[14\]\[31\] _1235_ _3396_ _3431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4632__S _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6716__A1 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6132__B _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7516__I0 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5690__C _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__S _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_78_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4750__I0 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4079__S _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6026__C _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5865__C _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__S _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5638__S _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6042__B _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5881__B _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5240_ _1856_ _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_121_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5171_ _1093_ memory\[30\]\[0\] _1819_ _1820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4122_ _1247_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4717__S _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4053_ net11 _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_69_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput3 address_i[2] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_79_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7812_ _0112_ clknet_leaf_129_clk_i memory\[29\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7743_ _0043_ clknet_leaf_182_clk_i memory\[19\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4955_ _1704_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4452__S _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3906_ memory\[19\]\[0\] _1093_ _1098_ _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7674_ _3836_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4886_ _1082_ memory\[25\]\[27\] _1660_ _1668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6625_ memory\[14\]\[28\] _3214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_89_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6556_ _1864_ memory\[6\]\[26\] _3147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_131_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5507_ memory\[16\]\[4\] memory\[17\]\[4\] _1911_ _2120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6487_ _2754_ _3078_ _2666_ _3079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8226_ _0526_ clknet_leaf_152_clk_i memory\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5438_ _2005_ _2007_ memory\[5\]\[2\] _2053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4732__I0 _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5369_ _1934_ _1984_ _1937_ _1985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8157_ _0457_ clknet_leaf_4_clk_i memory\[26\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8088_ _0388_ clknet_leaf_9_clk_i memory\[24\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7108_ memory\[31\]\[28\] _1229_ _3528_ _3537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5437__A1 _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7039_ memory\[13\]\[28\] _1229_ _3491_ _3500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_98_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4362__S _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7673__S _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_131_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5676__A1 _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4723__I0 _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__A2 _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_105_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6752__S _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5368__S _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4272__S _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4740_ _1076_ memory\[23\]\[24\] _1584_ _1589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4671_ _1551_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6410_ _2626_ memory\[19\]\[23\] _3003_ _2003_ _3004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_7390_ _1093_ memory\[0\]\[0\] _3686_ _3687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7583__S _3781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4071__I net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ _2515_ memory\[7\]\[21\] _2936_ _2517_ _2937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_clkbuf_leaf_101_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4962__I0 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6272_ _1094_ _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_40_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5667__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6927__S _3433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8011_ _0311_ clknet_leaf_45_clk_i memory\[22\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5223_ _1150_ memory\[30\]\[25\] _1841_ _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5154_ _1810_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4105_ net30 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6092__A1 _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5085_ _1076_ memory\[28\]\[24\] _1769_ _1774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4036_ _1188_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5786__B _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_26_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5987_ memory\[14\]\[14\] _2590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_94_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6395__A2 _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7726_ _0026_ clknet_leaf_89_clk_i memory\[19\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4938_ _1695_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4182__S _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4869_ _1056_ memory\[25\]\[19\] _1649_ _1659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7657_ memory\[6\]\[30\] net29 _3794_ _3828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7493__S _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6608_ _2803_ _1990_ memory\[25\]\[28\] _3197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4910__S _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7588_ _3791_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6539_ _3127_ _3129_ _2768_ _3130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_91_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5658__A1 _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8209_ _0509_ clknet_leaf_46_clk_i memory\[28\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6837__S _3383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5130__I0 _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5830__A1 _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6304__C _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3995__I1 _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4820__S _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_15_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4944__I0 _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6320__B _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6747__S _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7110__I1 _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5121__I0 _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6074__A1 _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5910_ _1861_ _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_88_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6890_ _3421_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5841_ _2160_ memory\[19\]\[11\] _2446_ _2075_ _2447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_88_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8560_ _0860_ clknet_leaf_96_clk_i memory\[3\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5772_ _1855_ _2355_ _2378_ _2379_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4723_ _1273_ memory\[23\]\[16\] _1573_ _1580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8491_ _0791_ clknet_leaf_84_clk_i memory\[11\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3986__I1 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7511_ _3750_ _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7442_ _1150_ memory\[0\]\[25\] _3708_ _3714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4654_ _1542_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5888__A1 _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4585_ _1505_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4935__I0 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_205_clk_i clknet_4_2_0_clk_i clknet_leaf_205_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7373_ _3677_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6324_ memory\[12\]\[21\] memory\[13\]\[21\] _2919_ _2920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6255_ _2803_ _2526_ memory\[25\]\[20\] _2852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_12_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5206_ _1133_ memory\[30\]\[17\] _1830_ _1838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6301__A2 _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6186_ _2784_ memory\[0\]\[18\] _2785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5137_ _1801_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5068_ _1273_ memory\[28\]\[16\] _1758_ _1765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input14_I data_i[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4019_ net31 _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_94_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3977__I1 _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7709_ _0009_ clknet_leaf_196_clk_i memory\[7\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8689_ _0989_ clknet_leaf_69_clk_i memory\[5\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5179__I0 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7168__I1 _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5963__C _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5879__A1 _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5270__I _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6366__I _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6056__A1 _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5103__I0 _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5803__A1 _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7398__S _3686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3968__I1 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4370_ _1390_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6295__A1 _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_191_clk_i clknet_4_3_0_clk_i clknet_leaf_191_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6040_ memory\[8\]\[15\] memory\[9\]\[15\] _2314_ _2642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_72_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input6_I data_i[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6047__A1 _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6209__C _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7991_ _0291_ clknet_leaf_41_clk_i memory\[21\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6942_ _1127_ memory\[16\]\[14\] _3444_ _3449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4725__S _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6873_ _3412_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_124_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6940__S _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5824_ _2380_ _2404_ _2429_ _2430_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_8612_ _0912_ clknet_leaf_144_clk_i memory\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5755_ _2362_ memory\[10\]\[9\] _2363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8543_ _0843_ clknet_leaf_168_clk_i memory\[8\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5783__C _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4706_ _1256_ memory\[23\]\[8\] _1562_ _1571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5686_ memory\[20\]\[8\] memory\[21\]\[8\] _1897_ _2295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_144_clk_i clknet_4_11_0_clk_i clknet_leaf_144_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_45_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8474_ _0774_ clknet_leaf_4_clk_i memory\[31\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7425_ _1133_ memory\[0\]\[17\] _3697_ _3705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4637_ _1533_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4908__I0 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5325__A3 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7356_ _3668_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4568_ _1496_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_9_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7287_ _1131_ memory\[3\]\[16\] _3625_ _3632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4499_ _1459_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6307_ _2574_ memory\[28\]\[21\] _2903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_159_clk_i clknet_4_10_0_clk_i clknet_leaf_159_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6286__A1 _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6238_ memory\[2\]\[19\] memory\[3\]\[19\] _2736_ _2836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6169_ _1915_ _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6119__C _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3895__I0 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6833__I0 _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5265__I _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6513__A2 _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_148_clk_i_I clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6277__B2 _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_200_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3870_ _1072_ memory\[7\]\[22\] _1066_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_61_clk_i clknet_4_7_0_clk_i clknet_leaf_61_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_73_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5540_ _2063_ memory\[29\]\[5\] _2151_ _1880_ _2152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4280__S _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5471_ _1930_ memory\[10\]\[3\] _2085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_54_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7210_ _3591_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7552__I1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4422_ _1418_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7591__S _3758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_76_clk_i clknet_4_6_0_clk_i clknet_leaf_76_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8190_ _0490_ clknet_leaf_15_clk_i memory\[27\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7141_ memory\[11\]\[11\] _1194_ _3553_ _3555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4353_ _1381_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_120_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7072_ _3518_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4284_ _1252_ memory\[17\]\[6\] _1336_ _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6268__A1 _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6023_ _2622_ _2294_ _2624_ _2250_ _2625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5778__C _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_14_clk_i clknet_4_1_0_clk_i clknet_leaf_14_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7974_ _0274_ clknet_leaf_161_clk_i memory\[21\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4455__S _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6925_ _1110_ memory\[16\]\[6\] _3433_ _3440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_85_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6440__A1 _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5243__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7240__I0 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6856_ _3403_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5794__B _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6787_ _1108_ memory\[9\]\[5\] _3361_ _3367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5807_ _1889_ _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_29_clk_i clknet_4_6_0_clk_i clknet_leaf_29_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6743__A2 _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3999_ _1161_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8526_ _0826_ clknet_leaf_98_clk_i memory\[8\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5738_ _1059_ _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_70_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4190__S _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7543__I1 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5669_ _2261_ _2266_ _2273_ _2278_ _1952_ _2279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_8457_ _0757_ clknet_leaf_127_clk_i memory\[31\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7408_ _1116_ memory\[0\]\[9\] _3686_ _3696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8388_ _0688_ clknet_leaf_141_clk_i memory\[16\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7339_ _3659_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_96_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7006__S _3480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6259__A1 _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6845__S _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6806__I0 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4365__S _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5688__C _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6431__A1 _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7676__S _3837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4293__I0 _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_74_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5196__S _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_109_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6734__A2 _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6498__B2 _3089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_118_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_56_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7298__I0 _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7470__I0 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6422__A1 _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4284__I0 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4971_ memory\[27\]\[2\] _1175_ _1711_ _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_127_Left_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7690_ _1127_ memory\[7\]\[14\] _3837_ _3845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3922_ _1109_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6490__S _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6710_ memory\[12\]\[30\] memory\[13\]\[30\] _2919_ _3297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3853_ net1 _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_74_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6641_ _2981_ memory\[7\]\[28\] _3229_ _2983_ _3230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_117_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _3159_ _3161_ _2757_ _3162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8311_ _0611_ clknet_leaf_18_clk_i net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5523_ _1238_ _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8242_ _0542_ clknet_leaf_83_clk_i memory\[2\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5454_ _1883_ _2067_ _1887_ _2068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_136_Left_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8173_ _0473_ clknet_leaf_56_clk_i memory\[27\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5385_ _1863_ _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4405_ _1408_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7289__I0 _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7124_ memory\[11\]\[3\] _1177_ _3542_ _3546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4336_ _1091_ memory\[17\]\[31\] _1335_ _1370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7055_ _3509_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4267_ _1333_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4511__I1 _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6006_ _2467_ _2605_ _2607_ _2608_ _2609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4198_ _1059_ _1295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XANTENNA__6661__A1 _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7957_ _0257_ clknet_leaf_35_clk_i memory\[20\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7888_ _0188_ clknet_leaf_70_clk_i memory\[18\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6908_ _3430_ _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7213__I0 _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6839_ _1160_ memory\[9\]\[30\] _3360_ _3394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_134_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6413__B _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7295__I _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4578__I1 _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5744__S _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8509_ _0809_ clknet_leaf_198_clk_i memory\[11\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6652__A1 _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7452__I0 _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4266__I0 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7204__I0 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4569__I1 _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5654__S _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5170_ _1818_ _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4121_ _1246_ memory\[15\]\[3\] _1240_ _1247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4052_ _1199_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6643__A1 _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 address_i[3] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6217__C _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7811_ _0111_ clknet_leaf_136_clk_i memory\[29\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7742_ _0042_ clknet_leaf_186_clk_i memory\[19\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4954_ _1082_ memory\[26\]\[27\] _1696_ _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3905_ _1097_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_52_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7673_ _1110_ memory\[7\]\[6\] _1087_ _3836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ _1667_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6624_ _3198_ _3203_ _3207_ _3212_ _2869_ _3213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5564__S _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6555_ memory\[4\]\[26\] _2934_ _3146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5506_ _1904_ memory\[19\]\[4\] _2118_ _2075_ _2119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8225_ _0525_ clknet_leaf_140_clk_i memory\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6486_ memory\[30\]\[25\] memory\[31\]\[25\] _1923_ _3078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5437_ _2049_ memory\[7\]\[2\] _2050_ _2051_ _2052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_clkbuf_leaf_22_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5368_ memory\[8\]\[1\] memory\[9\]\[1\] _1935_ _1984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8156_ _0456_ clknet_leaf_6_clk_i memory\[26\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4319_ _1361_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8087_ _0387_ clknet_leaf_10_clk_i memory\[24\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7107_ _3536_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4908__S _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5299_ _1915_ _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7682__I0 _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6634__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7038_ _3499_ _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6127__C _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4248__I0 _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7434__I0 _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4643__S _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5739__S _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4799__I1 _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5373__A1 _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4971__I1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5273__I _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4479__A3 _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4818__S _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7673__I0 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7425__I0 _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4239__I0 _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4553__S _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5649__S _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4670_ memory\[22\]\[24\] _1221_ _1546_ _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5892__B _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5364__B2 _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6340_ _2562_ memory\[6\]\[21\] _2936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_116_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6271_ _2865_ _2867_ _2768_ _2868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_11_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5667__A2 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8010_ _0310_ clknet_leaf_82_clk_i memory\[22\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5222_ _1846_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_196_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_135_Right_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5153_ _1148_ memory\[2\]\[24\] _1805_ _1810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4104_ _1234_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7104__S _3528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5084_ _1773_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4035_ memory\[12\]\[8\] _1187_ _1171_ _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4463__S _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5986_ _2573_ _2579_ _2583_ _2588_ _2403_ _2589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_75_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7725_ _0025_ clknet_leaf_101_clk_i memory\[19\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4937_ _1056_ memory\[26\]\[19\] _1685_ _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4868_ _1658_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7656_ _3827_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6147__A3 _2745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6607_ _2848_ memory\[27\]\[28\] _3195_ _2850_ _3196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_7_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5355__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4799_ memory\[24\]\[18\] _1208_ _1613_ _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4402__I0 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7587_ memory\[5\]\[29\] net27 _3781_ _3791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6410__C _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6538_ _1873_ _3128_ _2961_ _3129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6469_ _2884_ _3061_ _1913_ _3062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8208_ _0508_ clknet_leaf_46_clk_i memory\[28\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8139_ _0439_ clknet_leaf_45_clk_i memory\[26\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4638__S _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7014__S _3480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5821__I _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6607__A1 _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6138__B _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4469__I0 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6083__A2 _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6853__S _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4373__S _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7684__S _3837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5268__I _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5346__A1 _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5897__A2 _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__B _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4880__I0 _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5840_ _2208_ memory\[18\]\[11\] _2446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_88_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5771_ _2330_ net70 _2379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5585__A1 _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4722_ _1579_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8490_ _0790_ clknet_leaf_85_clk_i memory\[11\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7510_ _1150_ memory\[10\]\[25\] _3744_ _3750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7441_ _3713_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4653_ memory\[22\]\[16\] _1204_ _1535_ _1542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6511__B _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4584_ memory\[21\]\[16\] _1204_ _1498_ _1505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_77_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7372_ _1148_ memory\[4\]\[24\] _3672_ _3677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6938__S _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6323_ _1884_ _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5842__S _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6254_ _2848_ memory\[27\]\[20\] _2849_ _2850_ _2851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_40_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5205_ _1837_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ _1869_ _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5136_ _1273_ memory\[2\]\[16\] _1794_ _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_4_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5067_ _1764_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6673__S _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4018_ _1176_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_88_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7568__I _3758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5576__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5969_ _2337_ _2526_ memory\[25\]\[14\] _2572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_23_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4921__S _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7708_ _0008_ clknet_leaf_2_clk_i memory\[7\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8688_ _0988_ clknet_leaf_67_clk_i memory\[5\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5328__A1 _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7639_ memory\[6\]\[21\] net19 _3817_ _3819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_121_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5551__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6851__I1 _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7478__I _3721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5500__B _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6315__C _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_144_clk_i_I clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6331__B _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_113_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_69_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5461__I _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4278__S _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6295__A2 _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7589__S _3758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7990_ _0290_ clknet_leaf_42_clk_i memory\[21\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6941_ _3448_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4853__I0 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6506__B _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6872_ memory\[14\]\[13\] _1198_ _3408_ _3412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_124_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5823_ _2330_ net40 _2430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8611_ _0911_ clknet_leaf_152_clk_i memory\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5837__S _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8542_ _0842_ clknet_leaf_168_clk_i memory\[8\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5754_ _1869_ _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_57_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5685_ _1893_ _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4705_ _1570_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8473_ _0773_ clknet_leaf_16_clk_i memory\[31\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7424_ _3704_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4636_ memory\[22\]\[8\] _1187_ _1524_ _1533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7355_ _1131_ memory\[4\]\[16\] _3661_ _3668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5730__A1 _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6668__S _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4567_ memory\[21\]\[8\] _1187_ _1487_ _1496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6306_ _2798_ _2897_ _2900_ _2901_ _2902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_9_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7286_ _3631_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4498_ memory\[20\]\[8\] _1187_ _1450_ _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5371__I _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6237_ _2733_ memory\[1\]\[19\] _2834_ _2509_ _2835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4188__S _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6168_ _2629_ _2766_ _2495_ _2767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5119_ _1256_ memory\[2\]\[8\] _1783_ _1792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4916__S _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6099_ _2684_ _2689_ _2694_ _2699_ _2428_ _2700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5097__I0 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5797__B2 _2402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4844__I0 _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6135__C _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5549__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4651__S _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7010__I1 _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_70_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6277__A2 _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7077__I1 _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4826__S _1601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7202__S _3578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7001__I _3468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_204_clk_i clknet_4_2_0_clk_i clknet_leaf_204_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6045__C _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4561__S _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4063__I1 _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_219_clk_i clknet_4_0_0_clk_i clknet_leaf_219_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5960__A1 _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5470_ _2081_ _1921_ _2083_ _1927_ _2084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_112_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4421_ _1248_ memory\[1\]\[4\] _1413_ _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7140_ _3554_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4352_ _1248_ memory\[18\]\[4\] _1376_ _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7071_ memory\[31\]\[10\] _1191_ _3517_ _3518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4283_ _1342_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5191__I _1818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5405__B _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6287__I _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6022_ memory\[23\]\[15\] _2247_ _2623_ _2205_ _2624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7068__I1 _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4736__S _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5079__I0 _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7112__S _3505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5779__A1 _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7973_ _0273_ clknet_leaf_161_clk_i memory\[21\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6924_ _3439_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6440__A2 _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__S _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6855_ memory\[14\]\[5\] _1181_ _3397_ _3403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4054__I1 _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5806_ _2313_ _2412_ _2177_ _2413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6786_ _3366_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3998_ memory\[19\]\[30\] _1160_ _1097_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8525_ _0825_ clknet_leaf_98_clk_i memory\[8\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5737_ memory\[22\]\[9\] _2345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8456_ _0756_ clknet_leaf_123_clk_i memory\[31\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5668_ _1997_ _2274_ _2276_ _2277_ _2278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_7407_ _3695_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5703__A1 _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5599_ _2160_ memory\[19\]\[6\] _2209_ _2075_ _2210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4619_ _1523_ _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8387_ _0687_ clknet_leaf_138_clk_i memory\[16\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7338_ _1114_ memory\[4\]\[8\] _3650_ _3659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7269_ _3622_ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6197__I _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7456__A1 _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6861__S _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5985__B _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4045__I1 _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4381__S _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6195__A1 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_190_clk_i clknet_4_3_0_clk_i clknet_leaf_190_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_125_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5942__B2 _2545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7692__S _3837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5879__C _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6670__A2 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_143_clk_i clknet_4_11_0_clk_i clknet_leaf_143_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_25_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _1713_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3921_ memory\[19\]\[5\] _1108_ _1098_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6186__A1 _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3852_ _1057_ _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__5233__I0 _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_158_clk_i clknet_4_10_0_clk_i clknet_leaf_158_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6640_ _1864_ memory\[6\]\[28\] _3229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_39_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6571_ _2754_ _3160_ _1856_ _3161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5522_ memory\[2\]\[4\] memory\[3\]\[4\] _1992_ _2135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8310_ _0610_ clknet_leaf_18_clk_i net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4090__I net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8241_ _0541_ clknet_leaf_93_clk_i memory\[2\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5453_ memory\[30\]\[3\] memory\[31\]\[3\] _2066_ _2067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8172_ _0472_ clknet_leaf_55_clk_i memory\[27\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4404_ _1086_ memory\[18\]\[29\] _1398_ _1408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5384_ _1861_ _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6946__S _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4335_ _1369_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7123_ _3545_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6110__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7054_ memory\[31\]\[2\] _1175_ _3506_ _3509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4266_ _1089_ memory\[29\]\[30\] _1299_ _1333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6005_ _2472_ _2473_ memory\[5\]\[14\] _2608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4197_ _1293_ _1165_ _1094_ _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_38_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7956_ _0256_ clknet_leaf_35_clk_i memory\[20\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7887_ _0187_ clknet_leaf_89_clk_i memory\[18\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6907_ memory\[14\]\[30\] _1233_ _3396_ _3430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6838_ _3393_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5924__A1 _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_98_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8508_ _0808_ clknet_leaf_212_clk_i memory\[11\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6769_ _1927_ _3351_ _3353_ _3354_ _3355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_116_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8439_ _0739_ clknet_leaf_6_clk_i memory\[13\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6101__A1 _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_60_clk_i clknet_4_7_0_clk_i clknet_leaf_60_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_75_clk_i clknet_4_6_0_clk_i clknet_leaf_75_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_16_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6168__A1 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5000__S _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5215__I0 _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5915__A1 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6963__I0 _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_13_clk_i clknet_4_1_0_clk_i clknet_leaf_13_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6340__A1 _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_28_clk_i clknet_4_6_0_clk_i clknet_leaf_28_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4120_ net31 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4051_ memory\[12\]\[13\] _1198_ _1192_ _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4286__S _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput5 address_i[4] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7810_ _0110_ clknet_leaf_135_clk_i memory\[29\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7597__S _3795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5603__B1 _2207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7741_ _0041_ clknet_leaf_184_clk_i memory\[19\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_192_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4953_ _1703_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7672_ _3835_ _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3904_ _1096_ _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_46_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5206__I0 _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6623_ _3209_ _3211_ _1915_ _3212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4884_ _1080_ memory\[25\]\[26\] _1660_ _1667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6554_ _3142_ _3144_ _2887_ _3145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_27_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5505_ _1905_ memory\[18\]\[4\] _2118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6485_ _2000_ memory\[29\]\[25\] _3076_ _2855_ _3077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5436_ _1866_ _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8224_ _0524_ clknet_leaf_133_clk_i memory\[28\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5367_ _1929_ memory\[11\]\[1\] _1982_ _1932_ _1983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8155_ _0455_ clknet_leaf_6_clk_i memory\[26\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4318_ _1072_ memory\[17\]\[22\] _1358_ _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5298_ net4 _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8086_ _0386_ clknet_leaf_11_clk_i memory\[24\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7106_ memory\[31\]\[27\] _1227_ _3528_ _3536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input37_I data_i[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4249_ _1324_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7037_ memory\[13\]\[27\] _1227_ _3491_ _3499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6408__C _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4496__I1 _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6398__A1 _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7300__S _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7939_ _0239_ clknet_leaf_166_clk_i memory\[20\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7198__I0 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5982__C _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4184__I0 _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7370__I0 _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__S _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6389__A1 _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__I _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_64_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6936__I0 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6561__A1 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5364__A2 _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7361__I0 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6270_ _2629_ _2866_ _2495_ _2867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_139_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5221_ _1148_ memory\[30\]\[24\] _1841_ _1846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5152_ _1809_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4103_ memory\[12\]\[30\] _1233_ _1170_ _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5083_ _1074_ memory\[28\]\[23\] _1769_ _1773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4034_ net36 _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4744__S _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7120__S _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5985_ _2585_ _2587_ _2302_ _2588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7724_ _0024_ clknet_leaf_101_clk_i memory\[19\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4936_ _1694_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6927__I0 _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4867_ _1277_ memory\[25\]\[18\] _1649_ _1658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7655_ memory\[6\]\[29\] net27 _3817_ _3827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6606_ _2898_ memory\[26\]\[28\] _3195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_7_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7586_ _3790_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4798_ _1621_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6537_ memory\[16\]\[26\] memory\[17\]\[26\] _1885_ _3128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5374__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6304__A1 _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6468_ memory\[2\]\[24\] memory\[3\]\[24\] _2736_ _3061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8207_ _0507_ clknet_leaf_46_clk_i memory\[28\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4919__S _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6399_ _2798_ _2989_ _2991_ _2992_ _2993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5419_ memory\[12\]\[2\] memory\[13\]\[2\] _1978_ _2034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8138_ _0438_ clknet_leaf_177_clk_i memory\[26\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5323__B _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8069_ _0369_ clknet_leaf_155_clk_i memory\[24\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7655__I1 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5291__A1 _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6933__I _3432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4641__I1 _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_12_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6543__B2 _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5284__I _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7343__I0 _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_140_clk_i_I clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_65_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5770_ _2361_ _2367_ _2372_ _2377_ _1952_ _2378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_8_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4632__I1 _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4721_ _1271_ memory\[23\]\[15\] _1573_ _1579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_123_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4652_ _1541_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7440_ _1148_ memory\[0\]\[24\] _3708_ _3713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4396__I0 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput30 data_i[31] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4583_ _1504_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_77_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7371_ _3676_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7334__I0 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6322_ memory\[14\]\[21\] _2918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_122_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ _1060_ _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5204_ _1131_ memory\[30\]\[16\] _1830_ _1837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5922__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6239__B _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6184_ _2778_ _2782_ _2414_ _2783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5135_ _1800_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7637__I1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5066_ _1271_ memory\[28\]\[15\] _1758_ _1764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5797__C _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4320__I0 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4017_ memory\[12\]\[2\] _1175_ _1171_ _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5968_ _2382_ memory\[27\]\[14\] _2570_ _2384_ _2571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5576__A2 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6773__A1 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4919_ _1260_ memory\[26\]\[10\] _1685_ _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7707_ _0007_ clknet_leaf_208_clk_i memory\[7\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5899_ _2310_ memory\[11\]\[12\] _2503_ _2174_ _2504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8687_ _0987_ clknet_leaf_68_clk_i memory\[5\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6525__A1 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7638_ _3818_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7569_ memory\[5\]\[20\] net18 _3781_ _3782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4649__S _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4139__I0 _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7025__S _3491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7628__I1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6056__A3 _2656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4311__I0 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5264__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5279__I _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6516__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7316__I0 _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4559__S _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6940_ _1125_ memory\[16\]\[13\] _3444_ _3448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _3411_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_124_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5410__C _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5822_ _2409_ _2415_ _2422_ _2427_ _2428_ _2429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_8610_ _0910_ clknet_leaf_141_clk_i memory\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6755__A1 _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4093__I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__I1 _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5753_ _2356_ _1921_ _2359_ _2360_ _2361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_9_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8541_ _0841_ clknet_leaf_168_clk_i memory\[8\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4704_ _1254_ memory\[23\]\[7\] _1562_ _1570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5684_ memory\[22\]\[8\] _2293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8472_ _0772_ clknet_leaf_4_clk_i memory\[31\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5853__S _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7423_ _1131_ memory\[0\]\[16\] _3697_ _3704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4369__I0 _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4635_ _1532_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7354_ _3667_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4566_ _1495_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6305_ _2803_ _2526_ memory\[25\]\[21\] _2901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5730__A2 _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4469__S _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7285_ _1129_ memory\[3\]\[15\] _3625_ _3631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4497_ _1458_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6236_ _2784_ memory\[0\]\[19\] _2834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5494__A1 _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6167_ memory\[16\]\[18\] memory\[17\]\[18\] _2630_ _2766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5118_ _1791_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6098_ _2467_ _2695_ _2697_ _2698_ _2699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5601__B _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5049_ _1254_ memory\[28\]\[7\] _1747_ _1755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6746__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8739_ _1039_ clknet_leaf_120_clk_i memory\[7\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4731__I _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6859__S _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5990__C _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5021__I1 _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4379__S _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5562__I _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_13_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5485__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6594__S _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6326__C _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6737__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4842__S _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4420_ _1417_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_124_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4351_ _1380_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4282_ _1250_ memory\[17\]\[5\] _1336_ _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7070_ _3505_ _3517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_1_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6021_ memory\[20\]\[15\] memory\[21\]\[15\] _2346_ _2623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5476__A1 _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3921__S _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5779__A2 _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7972_ _0272_ clknet_leaf_161_clk_i memory\[21\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6923_ _1108_ memory\[16\]\[5\] _3433_ _3439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_85_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4826__I1 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5848__S _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4752__S _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6854_ _3402_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5805_ memory\[8\]\[10\] memory\[9\]\[10\] _2314_ _2412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6785_ _1106_ memory\[9\]\[4\] _3361_ _3366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3997_ net29 _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5400__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8524_ _0824_ clknet_leaf_97_clk_i memory\[8\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5736_ _2341_ _2343_ _2291_ _2344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5667_ _2005_ _2007_ memory\[5\]\[7\] _2277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8455_ _0755_ clknet_leaf_123_clk_i memory\[31\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7406_ _1114_ memory\[0\]\[8\] _3686_ _3695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4618_ _1522_ _1448_ _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_32_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5598_ _2208_ memory\[18\]\[6\] _2209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8386_ _0686_ clknet_leaf_137_clk_i memory\[16\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7337_ _3658_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_96_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4549_ _1485_ _1448_ _1486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__5382__I _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7268_ _1112_ memory\[3\]\[7\] _3614_ _3622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_187_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4927__S _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6219_ _2626_ memory\[19\]\[19\] _2816_ _2541_ _2817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7199_ _3585_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6427__B _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__S _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6719__A1 _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6589__S _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5292__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6388__I _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5458__B2 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7213__S _3589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4808__I1 _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4572__S _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3920_ net33 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_98_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A1 _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3851_ net3 _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_128_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4197__A1 _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6570_ memory\[30\]\[27\] memory\[31\]\[27\] _1923_ _3160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_4_Left_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5521_ _1987_ memory\[1\]\[4\] _2133_ _2043_ _2134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_80_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6981__I1 _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8240_ _0540_ clknet_leaf_96_clk_i memory\[2\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5452_ _1884_ _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_41_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8171_ _0471_ clknet_leaf_45_clk_i memory\[27\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5383_ memory\[4\]\[1\] _1998_ _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4744__I0 _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4403_ _1407_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5416__B _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4334_ _1089_ memory\[17\]\[30\] _1335_ _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7122_ memory\[11\]\[2\] _1175_ _3542_ _3545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7053_ _3508_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6004_ _2515_ memory\[7\]\[14\] _2606_ _2517_ _2607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4265_ _1332_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4196_ net3 _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5621__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7955_ _0255_ clknet_leaf_42_clk_i memory\[20\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4482__S _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7886_ _0186_ clknet_leaf_89_clk_i memory\[18\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6906_ _3429_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_108_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6837_ _1158_ memory\[9\]\[29\] _3383_ _3393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8507_ _0807_ clknet_leaf_215_clk_i memory\[11\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6768_ _1871_ _1934_ memory\[5\]\[31\] _3354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5719_ _1997_ _2324_ _2326_ _2327_ _2328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6699_ memory\[22\]\[30\] _3286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8438_ _0738_ clknet_leaf_5_clk_i memory\[13\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8369_ _0669_ clknet_leaf_67_clk_i memory\[14\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_203_clk_i clknet_4_2_0_clk_i clknet_leaf_203_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_130_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4657__S _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_9_clk_i clknet_4_1_0_clk_i clknet_leaf_9_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7033__S _3491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6157__B _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_218_clk_i clknet_4_0_0_clk_i clknet_leaf_218_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6872__S _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4392__S _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5287__I _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4567__S _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4050_ net10 _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6067__B _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5151__I0 _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5851__A1 _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 data_i[0] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5603__A1 _2196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_135_clk_i_I clknet_4_9_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7740_ _0040_ clknet_leaf_184_clk_i memory\[19\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4952_ _1080_ memory\[26\]\[26\] _1696_ _1703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7671_ _1108_ memory\[7\]\[5\] _1087_ _3835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3903_ _1062_ _1095_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4883_ _1666_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6622_ _1873_ _3210_ _2961_ _3211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5925__I _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6530__B _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6553_ _2884_ _3143_ _1913_ _3144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7118__S _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6484_ _2001_ memory\[28\]\[25\] _3076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_43_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5504_ _2114_ _1894_ _2116_ _1901_ _2117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__4717__I0 _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5435_ _2001_ memory\[6\]\[2\] _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8223_ _0523_ clknet_leaf_182_clk_i memory\[28\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6957__S _3455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5366_ _1930_ memory\[10\]\[1\] _1982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8154_ _0454_ clknet_leaf_5_clk_i memory\[26\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3940__I1 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5660__I _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8085_ _0385_ clknet_leaf_14_clk_i memory\[24\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4317_ _1360_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5297_ _1909_ _1912_ _1913_ _1914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4477__S _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7105_ _3535_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6095__A1 _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5142__I0 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4248_ _1070_ memory\[29\]\[21\] _1322_ _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7036_ _3498_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4179_ _1284_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6398__A2 _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_67_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7938_ _0238_ clknet_leaf_166_clk_i memory\[20\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4940__S _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7869_ _0169_ clknet_leaf_186_clk_i memory\[17\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4956__I0 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4708__I0 _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_142_clk_i clknet_4_11_0_clk_i clknet_leaf_142_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_76_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7122__I1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_157_clk_i clknet_4_10_0_clk_i clknet_leaf_157_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7698__S _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_85_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5011__S _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3998__I1 _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_64_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6561__A2 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6777__S _3361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ _1845_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_61_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4297__S _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5151_ _1146_ memory\[2\]\[23\] _1805_ _1809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5124__I0 _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6077__A1 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5082_ _1772_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4102_ net29 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6509__C _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5824__A1 _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4033_ _1186_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4096__I net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6017__S _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5984_ _2163_ _2586_ _2495_ _2587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7723_ _0023_ clknet_leaf_102_clk_i memory\[19\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3989__I1 _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4935_ _1277_ memory\[26\]\[18\] _1685_ _1694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4866_ _1657_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7654_ _3826_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4797_ memory\[24\]\[17\] _1206_ _1613_ _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6605_ memory\[24\]\[28\] _2799_ _3194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7585_ memory\[5\]\[28\] net26 _3781_ _3790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6536_ _1876_ memory\[19\]\[26\] _3126_ _2003_ _3127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_43_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6467_ _2733_ memory\[1\]\[24\] _3059_ _2975_ _3060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8206_ _0506_ clknet_leaf_73_clk_i memory\[28\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_74_clk_i clknet_4_6_0_clk_i clknet_leaf_74_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6398_ _2803_ _1990_ memory\[25\]\[23\] _2992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5418_ memory\[14\]\[2\] _2033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5349_ _1883_ _1964_ _1887_ _1965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8137_ _0437_ clknet_leaf_177_clk_i memory\[26\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5115__I0 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7104__I1 _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_89_clk_i clknet_4_13_0_clk_i clknet_leaf_89_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8068_ _0368_ clknet_leaf_163_clk_i memory\[24\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4935__S _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7019_ _3489_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_12_clk_i clknet_4_1_0_clk_i clknet_leaf_12_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6154__C _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4670__S _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4929__I0 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5565__I _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6170__B _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_27_clk_i clknet_4_6_0_clk_i clknet_leaf_27_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_80_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7591__I1 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6543__A2 _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6059__A1 _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5006__S _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5806__A1 _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7221__S _3589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6231__A1 _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4580__S _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4720_ _1578_ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6909__I1 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4651_ memory\[22\]\[15\] _1202_ _1535_ _1541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput31 data_i[3] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6534__A2 _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput20 data_i[22] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4582_ memory\[21\]\[15\] _1202_ _1498_ _1504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_77_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7370_ _1146_ memory\[4\]\[23\] _3672_ _3676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_123_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3924__S _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6321_ _2902_ _2907_ _2911_ _2916_ _2869_ _2917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_40_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6252_ _2432_ memory\[26\]\[20\] _2849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5203_ _1836_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_90_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6183_ _2779_ _2781_ _2643_ _2782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5134_ _1271_ memory\[2\]\[15\] _1794_ _1800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _1763_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4016_ net28 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_88_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7270__I0 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ _2432_ memory\[26\]\[14\] _2570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8755_ _1055_ clknet_leaf_83_clk_i memory\[7\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6773__A2 _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8686_ _0986_ clknet_leaf_68_clk_i memory\[5\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4918_ _1673_ _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_47_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4490__S _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7706_ _0006_ clknet_leaf_211_clk_i memory\[7\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_133_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5898_ _2362_ memory\[10\]\[12\] _2503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_118_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6702__C _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7637_ memory\[6\]\[20\] net18 _3817_ _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4849_ _1648_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5385__I _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7573__I1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7568_ _3758_ _3781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6519_ _2796_ net56 _3111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7499_ _3721_ _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6210__S _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7306__S _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6289__A1 _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5334__B _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3898__I0 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7041__S _3491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6461__A1 _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6880__S _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5509__B _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7564__I1 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6516__A2 _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6120__S _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6059__C _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6827__I0 _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6452__A1 _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ memory\[14\]\[12\] _1196_ _3408_ _3411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6204__A1 _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5821_ _1063_ _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5963__B1 _2560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5752_ _1058_ _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_8540_ _0840_ clknet_leaf_206_clk_i memory\[8\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4703_ _1569_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5683_ _2287_ _2290_ _2291_ _2292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8471_ _0771_ clknet_leaf_17_clk_i memory\[31\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7422_ _3703_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4634_ memory\[22\]\[7\] _1185_ _1524_ _1532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7353_ _1129_ memory\[4\]\[15\] _3661_ _3667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_102_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4565_ memory\[21\]\[7\] _1185_ _1487_ _1495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6304_ _2848_ memory\[27\]\[21\] _2899_ _2850_ _2900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7126__S _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7284_ _3630_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4496_ memory\[20\]\[7\] _1185_ _1450_ _1458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6235_ _2830_ _2832_ _2414_ _2833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6965__S _3455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_31_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6166_ _2626_ memory\[19\]\[18\] _2764_ _2541_ _2765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6691__A1 _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6097_ _2472_ _2473_ memory\[5\]\[16\] _2698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5117_ _1254_ memory\[2\]\[7\] _1783_ _1791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7491__I0 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5048_ _1754_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6443__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input12_I data_i[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_183_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_40_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8738_ _1038_ clknet_leaf_144_clk_i memory\[7\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6999_ memory\[13\]\[9\] _1189_ _3469_ _3479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8669_ _0969_ clknet_leaf_199_clk_i memory\[10\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4780__I1 _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4532__I1 _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5485__A2 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6682__A1 _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6607__C _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7234__I0 _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6623__B _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4599__I1 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5954__S _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7537__I1 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4220__I0 _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4350_ _1246_ memory\[18\]\[3\] _1376_ _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6785__S _3361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4281_ _1341_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6020_ memory\[22\]\[15\] _2622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input4_I address_i[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6425__A1 _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7971_ _0271_ clknet_leaf_166_clk_i memory\[21\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5421__C _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6922_ _3438_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7225__I0 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6853_ memory\[14\]\[4\] _1179_ _3397_ _3402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5804_ _2310_ memory\[11\]\[10\] _2410_ _2174_ _2411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_77_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5928__I _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6784_ _3365_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3996_ _1159_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5400__A2 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8523_ _0823_ clknet_leaf_89_clk_i memory\[8\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5735_ _2288_ _2342_ _2200_ _2343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5666_ _2049_ memory\[7\]\[7\] _2275_ _2051_ _2276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8454_ _0754_ clknet_leaf_122_clk_i memory\[31\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7405_ _3694_ _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4617_ net38 _1372_ _1522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_45_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5597_ _1863_ _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_8385_ _0685_ clknet_leaf_137_clk_i memory\[16\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7336_ _1112_ memory\[4\]\[7\] _3650_ _3658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_96_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4548_ net38 _1296_ _1485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__4762__I1 _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7267_ _3621_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4479_ _1057_ _1165_ _1063_ _1448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_96_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6218_ _2674_ memory\[18\]\[19\] _2816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6664__A1 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5612__B _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7198_ _1110_ memory\[8\]\[6\] _3578_ _3585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6149_ _2432_ memory\[26\]\[18\] _2748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7464__I0 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4278__I0 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4450__I0 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5506__C _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4505__I1 _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6655__A1 _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5458__A2 _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6407__B2 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5949__S _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4853__S _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7207__I0 _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6072__C _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3850_ net16 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_46_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5520_ _1988_ memory\[0\]\[4\] _2133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__I1 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5451_ _2063_ memory\[29\]\[3\] _2064_ _1880_ _2065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_131_clk_i_I clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5382_ _1858_ _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4402_ _1084_ memory\[18\]\[28\] _1398_ _1407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8170_ _0470_ clknet_leaf_177_clk_i memory\[27\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7121_ _3544_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4333_ _1368_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4099__I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7694__I0 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7404__S _3686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7052_ memory\[31\]\[1\] _1173_ _3506_ _3508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4264_ _1086_ memory\[29\]\[29\] _1322_ _1332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6003_ _2562_ memory\[6\]\[14\] _2606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5432__B _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_105_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_4_14_0_clk_i clknet_0_clk_i clknet_4_14_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4195_ _1292_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7446__I0 _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7954_ _0254_ clknet_leaf_44_clk_i memory\[20\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5621__A2 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6905_ memory\[14\]\[29\] _1231_ _3419_ _3429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7885_ _0185_ clknet_leaf_101_clk_i memory\[18\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_56_clk_i_I clknet_4_5_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6836_ _3392_ _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_114_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6767_ _2981_ memory\[7\]\[31\] _3352_ _2983_ _3353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_9_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5718_ _2005_ _2007_ memory\[5\]\[8\] _2327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_98_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8506_ _0806_ clknet_leaf_212_clk_i memory\[11\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3979_ net22 _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_116_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6698_ _3282_ _3284_ _1889_ _3285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4983__I1 _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5649_ memory\[12\]\[7\] memory\[13\]\[7\] _1978_ _2259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8437_ _0737_ clknet_leaf_191_clk_i memory\[13\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8368_ _0668_ clknet_leaf_64_clk_i memory\[14\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5688__A2 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7319_ _3648_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_123_Left_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8299_ _0599_ clknet_leaf_72_clk_i net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7314__S _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6637__A1 _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_130_Right_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_132_Left_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4423__I0 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6620__C _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__S _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4848__S _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7676__I0 _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 data_i[10] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4951_ _1702_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7670_ _3834_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3902_ net3 net4 _1094_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_4882_ _1078_ memory\[25\]\[25\] _1660_ _1666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6621_ memory\[16\]\[28\] memory\[17\]\[28\] _1885_ _3210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5367__A1 _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3927__S _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6552_ memory\[2\]\[26\] memory\[3\]\[26\] _2736_ _3143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6483_ _2798_ _3071_ _3073_ _3074_ _3075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5503_ memory\[23\]\[4\] _1896_ _2115_ _1899_ _2116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_5434_ _1861_ _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8222_ _0522_ clknet_leaf_22_clk_i memory\[28\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4342__A2 _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8153_ _0453_ clknet_leaf_9_clk_i memory\[26\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7134__S _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7667__I0 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6619__A1 _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7104_ memory\[31\]\[26\] _1225_ _3528_ _3535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5365_ _1977_ _1921_ _1980_ _1927_ _1981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8084_ _0384_ clknet_leaf_35_clk_i memory\[24\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4316_ _1070_ memory\[17\]\[21\] _1358_ _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5296_ _1238_ _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_10_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4247_ _1323_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6973__S _3455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7035_ memory\[13\]\[26\] _1225_ _3491_ _3498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7419__I0 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4178_ _1074_ memory\[15\]\[23\] _1280_ _1284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7937_ _0237_ clknet_leaf_167_clk_i memory\[20\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4292__I _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7868_ _0168_ clknet_leaf_185_clk_i memory\[17\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5358__A1 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6819_ _1139_ memory\[9\]\[20\] _3383_ _3384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_102_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6721__B _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7799_ _0099_ clknet_leaf_220_clk_i memory\[15\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__S _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5530__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6168__B _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4892__I0 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5298__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5349__A1 _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7219__S _3589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6010__A2 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4578__S _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5521__A1 _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6078__B _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5150_ _1808_ _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6793__S _3361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5081_ _1072_ memory\[28\]\[22\] _1769_ _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4101_ _1232_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6872__I1 _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4032_ memory\[12\]\[7\] _1185_ _1171_ _1186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5202__S _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5983_ memory\[16\]\[14\] memory\[17\]\[14\] _2164_ _2586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4934_ _1693_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7722_ _0022_ clknet_leaf_86_clk_i memory\[19\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_202_clk_i clknet_4_2_0_clk_i clknet_leaf_202_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_118_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4865_ _1275_ memory\[25\]\[17\] _1649_ _1657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7653_ memory\[6\]\[28\] net26 _3817_ _3826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5060__I0 _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ _1620_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_8_clk_i clknet_4_1_0_clk_i clknet_leaf_8_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7584_ _3789_ _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6604_ _2846_ _3172_ _3192_ _3193_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_132_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5760__A1 _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6535_ _1877_ memory\[18\]\[26\] _3126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_7_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_217_clk_i clknet_4_0_0_clk_i clknet_leaf_217_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8205_ _0505_ clknet_leaf_71_clk_i memory\[28\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6466_ _2784_ memory\[0\]\[24\] _3059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6397_ _2848_ memory\[27\]\[23\] _2990_ _2850_ _2991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5417_ _2016_ _2021_ _2025_ _2031_ _1918_ _2032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__4488__S _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5348_ memory\[30\]\[1\] memory\[31\]\[1\] _1885_ _1964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8136_ _0436_ clknet_leaf_139_clk_i memory\[26\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8067_ _0367_ clknet_leaf_164_clk_i memory\[24\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7018_ memory\[13\]\[18\] _1208_ _3480_ _3489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5279_ _1895_ _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4874__I0 _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6863__I1 _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6716__B _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5579__A1 _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7039__S _3491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5051__I0 _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6878__S _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5751__B2 _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4398__S _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__B2 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_178_clk_i_I clknet_4_9_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5514__C _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7502__S _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4865__I0 _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4861__S _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4650_ _1540_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7031__I1 _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput10 data_i[13] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5742__A1 _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput21 data_i[23] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4581_ _1503_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput32 data_i[4] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6320_ _2913_ _2915_ _2768_ _2916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_52_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6251_ _1295_ _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_58_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5202_ _1129_ memory\[30\]\[15\] _1830_ _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_110_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6182_ memory\[8\]\[18\] memory\[9\]\[18\] _2780_ _2781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5133_ _1799_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7098__I1 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3940__S _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5064_ _1269_ memory\[28\]\[14\] _1758_ _1763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6845__I1 _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4015_ _1174_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_141_clk_i clknet_4_11_0_clk_i clknet_leaf_141_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_118_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ memory\[24\]\[14\] _2333_ _2569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8754_ _1054_ clknet_leaf_76_clk_i memory\[7\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5897_ _2499_ _2406_ _2501_ _2360_ _2502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_8685_ _0985_ clknet_leaf_92_clk_i memory\[5\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5981__A1 _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6271__B _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4917_ _1684_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7705_ _0005_ clknet_leaf_210_clk_i memory\[7\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4848_ _1258_ memory\[25\]\[9\] _1638_ _1648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_51_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_156_clk_i clknet_4_10_0_clk_i clknet_leaf_156_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7636_ _3794_ _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_133_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5733__A1 _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7567_ _3780_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6781__I0 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ _1611_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7498_ _3743_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6518_ _3094_ _3099_ _3104_ _3109_ _2894_ _3110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6449_ memory\[23\]\[24\] _2713_ _3041_ _2671_ _3042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6289__A2 _2885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4011__S _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5107__S _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7089__I1 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8119_ _0419_ clknet_leaf_10_clk_i memory\[25\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7322__S _3650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4946__S _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6446__B _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5350__B _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_109_clk_i clknet_4_15_0_clk_i clknet_leaf_109_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5972__A1 _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5525__B _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6200__I _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5017__S _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_72_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7232__S _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4838__I0 _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6075__C _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5820_ _1997_ _2423_ _2425_ _2426_ _2427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xclkbuf_leaf_73_clk_i clknet_4_6_0_clk_i clknet_leaf_73_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4066__I1 _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5751_ memory\[15\]\[9\] _2357_ _2358_ _2307_ _2359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__7004__I1 _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8470_ _0770_ clknet_leaf_17_clk_i memory\[31\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4702_ _1252_ memory\[23\]\[6\] _1562_ _1569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7421_ _1129_ memory\[0\]\[15\] _3697_ _3703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5682_ _1889_ _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_60_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_88_clk_i clknet_4_12_0_clk_i clknet_leaf_88_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_71_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4633_ _1531_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7352_ _3666_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4564_ _1494_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7283_ _1127_ memory\[3\]\[14\] _3625_ _3630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6303_ _2898_ memory\[26\]\[21\] _2899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_12_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7206__I _3577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6234_ _2779_ _2831_ _2643_ _2832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_11_clk_i clknet_4_1_0_clk_i clknet_leaf_11_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4495_ _1457_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6165_ _2674_ memory\[18\]\[18\] _2764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4766__S _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6096_ _2515_ memory\[7\]\[16\] _2696_ _2517_ _2697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5116_ _1790_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_26_clk_i clknet_4_3_0_clk_i clknet_leaf_26_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5047_ _1252_ memory\[28\]\[6\] _1747_ _1754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6981__S _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4057__I1 _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_126_clk_i_I clknet_4_14_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6998_ _3478_ _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_137_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5949_ memory\[8\]\[13\] memory\[9\]\[13\] _2314_ _2553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8737_ _1037_ clknet_leaf_145_clk_i memory\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8668_ _0968_ clknet_leaf_212_clk_i memory\[10\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_133_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7619_ _3808_ _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8599_ _0899_ clknet_leaf_209_clk_i memory\[4\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_133_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6131__A1 _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4676__S _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7052__S _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6891__S _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4048__I1 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6198__A1 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5945__B2 _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4280_ _1248_ memory\[17\]\[4\] _1336_ _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4586__S _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6865__I _3396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4385__I _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7970_ _0270_ clknet_leaf_166_clk_i memory\[21\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6921_ _1106_ memory\[16\]\[4\] _3433_ _3438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6189__A1 _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6852_ _3401_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5803_ _2362_ memory\[10\]\[10\] _2410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5210__S _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5936__A1 _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8522_ _0822_ clknet_leaf_88_clk_i memory\[8\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6783_ _1104_ memory\[9\]\[3\] _3361_ _3365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3995_ memory\[19\]\[29\] _1158_ _1140_ _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_33_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5734_ memory\[30\]\[9\] memory\[31\]\[9\] _2066_ _2342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5665_ _2096_ memory\[6\]\[7\] _2275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8453_ _0753_ clknet_leaf_120_clk_i memory\[31\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_10_0_clk_i clknet_0_clk_i clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7404_ _1112_ memory\[0\]\[7\] _3686_ _3694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4616_ _1521_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8384_ _0684_ clknet_leaf_173_clk_i memory\[14\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7335_ _3657_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6361__B2 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5596_ _2203_ _1894_ _2206_ _1901_ _2207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__5880__S _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4547_ _1484_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_52_clk_i_I clknet_4_5_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7266_ _1110_ memory\[3\]\[6\] _3614_ _3621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4478_ _1447_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7197_ _3584_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6217_ _2811_ _2760_ _2814_ _2716_ _2815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4496__S _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6148_ memory\[24\]\[18\] _2333_ _2747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6708__C _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6079_ _2662_ _2668_ _2673_ _2679_ _2403_ _2680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_67_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6443__C _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5227__I0 _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5927__A1 _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6975__I0 _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6352__A1 _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6104__A1 _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6618__C _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6407__A2 _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7510__S _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5918__A1 _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4197__A3 _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_80_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5450_ _1877_ memory\[28\]\[3\] _2064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4401_ _1406_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5381_ _1058_ _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7120_ memory\[11\]\[1\] _1173_ _3542_ _3544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4332_ _1086_ memory\[17\]\[29\] _1358_ _1368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5713__B _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7051_ _3507_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4263_ _1331_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6002_ memory\[4\]\[14\] _2468_ _2605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4194_ _1091_ memory\[15\]\[31\] _1239_ _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7953_ _0253_ clknet_leaf_50_clk_i memory\[20\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6904_ _3428_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7884_ _0184_ clknet_leaf_101_clk_i memory\[18\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4680__I1 _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6957__I0 _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6835_ _1156_ memory\[9\]\[28\] _3383_ _3392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3978_ _1147_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6766_ _1864_ memory\[6\]\[31\] _3352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_128_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5717_ _2049_ memory\[7\]\[8\] _2325_ _2051_ _2326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_98_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6582__B2 _3171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8505_ _0805_ clknet_leaf_212_clk_i memory\[11\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6697_ _1932_ _3283_ _1856_ _3284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8436_ _0736_ clknet_leaf_28_clk_i memory\[13\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5648_ memory\[14\]\[7\] _2258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5607__C _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7382__I0 _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8367_ _0667_ clknet_leaf_66_clk_i memory\[14\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5579_ _1954_ net66 _2191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4896__A1 _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8298_ _0598_ clknet_leaf_127_clk_i net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7318_ _1162_ memory\[3\]\[31\] _3613_ _3648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7249_ _3611_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5115__S _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7330__S _3650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4954__S _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6454__B _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6948__I0 _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6325__B2 _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6628__A2 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5025__S _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 data_i[11] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7240__S _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6083__C _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4662__I1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4950_ _1078_ memory\[26\]\[25\] _1696_ _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3901_ _1063_ _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_4881_ _1665_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6620_ _1876_ memory\[19\]\[28\] _3208_ _2003_ _3209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_46_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6564__A1 _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5708__B _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6551_ _2733_ memory\[1\]\[26\] _3141_ _2975_ _3142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5502_ memory\[20\]\[4\] memory\[21\]\[4\] _1897_ _2115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6316__A1 _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6482_ _2803_ _1990_ memory\[25\]\[25\] _3074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7364__I0 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5433_ memory\[4\]\[2\] _1998_ _2048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8221_ _0521_ clknet_leaf_15_clk_i memory\[28\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4178__I0 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7415__S _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3943__S _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8152_ _0452_ clknet_leaf_10_clk_i memory\[26\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5364_ memory\[15\]\[1\] _1922_ _1979_ _1925_ _1980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4315_ _1359_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6539__B _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7103_ _3534_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8083_ _0383_ clknet_leaf_42_clk_i memory\[24\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5295_ memory\[16\]\[0\] memory\[17\]\[0\] _1911_ _1912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4246_ _1068_ memory\[29\]\[20\] _1322_ _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7034_ _3497_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4350__I0 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4177_ _1283_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4774__S _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4653__I1 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7936_ _0236_ clknet_leaf_179_clk_i memory\[1\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7867_ _0167_ clknet_leaf_188_clk_i memory\[17\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _3360_ _3383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_135_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7798_ _0098_ clknet_leaf_220_clk_i memory\[15\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6749_ _3332_ _3334_ _1915_ _3335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7355__I0 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6307__A1 _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4014__S _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4169__I0 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8419_ _0719_ clknet_leaf_156_clk_i memory\[13\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4684__S _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7060__S _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6184__B _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_174_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6546__A1 _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4859__S _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7649__I1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_99_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5080_ _1771_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4100_ memory\[12\]\[29\] _1231_ _1213_ _1232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5824__A3 _2429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4031_ net35 _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4332__I0 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5982_ _2160_ memory\[19\]\[14\] _2584_ _2541_ _2585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4933_ _1275_ memory\[26\]\[17\] _1685_ _1693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7721_ _0021_ clknet_leaf_125_clk_i memory\[19\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4864_ _1656_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7652_ _3825_ _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4795_ memory\[24\]\[16\] _1204_ _1613_ _1620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7583_ memory\[5\]\[27\] net25 _3781_ _3789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6603_ _2796_ net58 _3193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6113__I _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6534_ _3122_ _2760_ _3124_ _2716_ _3125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6465_ _3055_ _3057_ _2880_ _3058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7145__S _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8204_ _0504_ clknet_leaf_57_clk_i memory\[28\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5416_ _2027_ _2030_ _1916_ _2031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6396_ _2898_ memory\[26\]\[23\] _2990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_101_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5347_ _1876_ memory\[29\]\[1\] _1962_ _1880_ _1963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8135_ _0435_ clknet_leaf_139_clk_i memory\[26\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5278_ _1061_ _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8066_ _0366_ clknet_leaf_175_clk_i memory\[24\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5901__B _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input35_I data_i[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4229_ _1265_ memory\[29\]\[12\] _1311_ _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7017_ _3488_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5620__C _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7919_ _0219_ clknet_leaf_100_clk_i memory\[1\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4626__I1 _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7328__I0 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5751__A2 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5862__I _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5503__A2 _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4314__I0 _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7500__I0 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5102__I _1782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6767__A1 _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5990__A2 _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6519__A1 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 data_i[14] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4580_ memory\[21\]\[14\] _1200_ _1498_ _1503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput22 data_i[24] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput33 data_i[5] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6250_ memory\[24\]\[20\] _2799_ _2847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5201_ _1835_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6181_ _1910_ _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5132_ _1269_ memory\[2\]\[14\] _1794_ _1799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4305__I0 _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5258__A1 _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5063_ _1762_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6536__C _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5213__S _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6309__S _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4014_ memory\[12\]\[1\] _1173_ _1171_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5440__C _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6758__A1 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5965_ _2380_ _2546_ _2567_ _2568_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_8753_ _1053_ clknet_leaf_69_clk_i memory\[7\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5896_ memory\[15\]\[12\] _2357_ _2500_ _2307_ _2501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_118_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8684_ _0984_ clknet_leaf_92_clk_i memory\[5\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4916_ _1258_ memory\[26\]\[9\] _1674_ _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7704_ _0004_ clknet_leaf_2_clk_i memory\[7\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7635_ _3816_ _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4847_ _1647_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7566_ memory\[5\]\[19\] net16 _3770_ _3780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4778_ memory\[24\]\[8\] _1187_ _1602_ _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5682__I _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7497_ _1137_ memory\[10\]\[19\] _3733_ _3743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6517_ _2933_ _3105_ _3107_ _3108_ _3109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6448_ memory\[20\]\[24\] memory\[21\]\[24\] _2812_ _3041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_122_clk_i_I clknet_4_14_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5497__A1 _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6379_ _2784_ memory\[0\]\[22\] _2974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7603__S _3795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8118_ _0418_ clknet_leaf_11_clk_i memory\[25\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8049_ _0349_ clknet_leaf_50_clk_i memory\[23\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4962__S _1673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4761__I _1601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_47_clk_i_I clknet_4_5_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6889__S _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5793__S _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5806__B _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5488__A1 _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_201_clk_i clknet_4_2_0_clk_i clknet_leaf_201_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_72_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6637__B _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_7_clk_i clknet_4_1_0_clk_i clknet_leaf_7_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_89_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_216_clk_i clknet_4_0_0_clk_i clknet_leaf_216_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4872__S _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5412__A1 _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5750_ memory\[12\]\[9\] memory\[13\]\[9\] _1978_ _2358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5681_ _2288_ _2289_ _2200_ _2290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4701_ _1568_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7420_ _3702_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5015__I1 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4632_ memory\[22\]\[6\] _1183_ _1524_ _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5715__A2 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7351_ _1127_ memory\[4\]\[14\] _3661_ _3666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5208__S _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4563_ memory\[21\]\[6\] _1183_ _1487_ _1494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7282_ _3629_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6302_ _1910_ _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4112__S _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4494_ memory\[20\]\[6\] _1183_ _1450_ _1457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6233_ memory\[8\]\[19\] memory\[9\]\[19\] _2780_ _2831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5479__A1 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7423__S _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6140__A2 _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6164_ _2759_ _2760_ _2762_ _2716_ _2763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_6095_ _2562_ memory\[6\]\[16\] _2696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5115_ _1252_ memory\[2\]\[6\] _1783_ _1790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5046_ _1753_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6266__C _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5403__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6282__B _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6997_ memory\[13\]\[8\] _1187_ _3469_ _3478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5948_ _2310_ memory\[11\]\[13\] _2551_ _2174_ _2552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_48_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8736_ _1036_ clknet_leaf_179_clk_i memory\[6\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5879_ _2063_ memory\[29\]\[12\] _2483_ _2389_ _2484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5006__I1 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8667_ _0967_ clknet_leaf_215_clk_i memory\[10\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7618_ memory\[6\]\[11\] net8 _3806_ _3808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_106_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8598_ _0898_ clknet_leaf_193_clk_i memory\[4\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7549_ _3771_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3861__S _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6176__C _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5788__S _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5642__A1 _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4692__S _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6198__A2 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5945__A2 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6993__I1 _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7508__S _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_140_clk_i clknet_4_11_0_clk_i clknet_leaf_140_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4867__S _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7170__I1 _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5181__I0 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6367__B _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5881__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5271__B _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_155_clk_i clknet_4_10_0_clk_i clknet_leaf_155_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6920_ _3437_ _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6851_ memory\[14\]\[3\] _1177_ _3397_ _3401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5802_ _2405_ _2406_ _2408_ _2360_ _2409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_71_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8521_ _0821_ clknet_leaf_102_clk_i memory\[8\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6782_ _3364_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3994_ net27 _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_33_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3946__S _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5733_ _2063_ memory\[29\]\[9\] _2340_ _1880_ _2341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_72_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5664_ memory\[4\]\[7\] _1998_ _2274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8452_ _0752_ clknet_leaf_143_clk_i memory\[31\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7403_ _3693_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4615_ memory\[21\]\[31\] _1235_ _1486_ _1521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8383_ _0683_ clknet_leaf_172_clk_i memory\[14\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5595_ memory\[23\]\[6\] _1896_ _2204_ _2205_ _2206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_130_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7334_ _1110_ memory\[4\]\[6\] _3650_ _3657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_108_clk_i clknet_4_15_0_clk_i clknet_leaf_108_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6361__A2 _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4546_ memory\[20\]\[31\] _1235_ _1449_ _1484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_96_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7153__S _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7265_ _3620_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4477_ _1091_ memory\[1\]\[31\] _1412_ _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7196_ _1108_ memory\[8\]\[5\] _3578_ _3584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6216_ memory\[23\]\[19\] _2713_ _2813_ _2671_ _2814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5872__A1 _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6147_ _2380_ _2723_ _2745_ _2746_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6078_ _2676_ _2678_ _2302_ _2679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5624__A1 _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5029_ memory\[27\]\[30\] _1233_ _1710_ _1744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4017__S _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8719_ _1019_ clknet_leaf_69_clk_i memory\[6\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7328__S _3650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6740__B _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4738__I0 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6352__A2 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3961__I1 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_72_clk_i clknet_4_7_0_clk_i clknet_leaf_72_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5163__I0 _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4910__I0 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_87_clk_i clknet_4_12_0_clk_i clknet_leaf_87_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_25_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_10_clk_i clknet_4_1_0_clk_i clknet_leaf_10_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_73_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7238__S _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4729__I0 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_25_clk_i clknet_4_3_0_clk_i clknet_leaf_25_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_112_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4400_ _1082_ memory\[18\]\[27\] _1398_ _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5380_ _1991_ _1995_ _1950_ _1996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7143__I1 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3952__I1 _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4597__S _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4331_ _1367_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7050_ memory\[31\]\[0\] _1164_ _3506_ _3507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4262_ _1084_ memory\[29\]\[28\] _1322_ _1331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6646__A3 _3233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_169_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5854__A1 _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6001_ _2600_ _2603_ _2421_ _2604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4193_ _1291_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7952_ _0252_ clknet_leaf_51_clk_i memory\[20\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5221__S _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5606__B2 _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6544__C _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6903_ memory\[14\]\[28\] _1229_ _3419_ _3428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7883_ _0183_ clknet_leaf_101_clk_i memory\[18\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6116__I _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5909__A2 _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6834_ _3391_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3977_ memory\[19\]\[23\] _1146_ _1140_ _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6765_ memory\[4\]\[31\] _1859_ _3351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5716_ _2096_ memory\[6\]\[8\] _2325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_98_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8504_ _0804_ clknet_leaf_211_clk_i memory\[11\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_98_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8435_ _0735_ clknet_leaf_75_clk_i memory\[13\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6696_ memory\[30\]\[30\] memory\[31\]\[30\] _1923_ _3283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6987__S _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5647_ _2240_ _2245_ _2251_ _2256_ _1918_ _2257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8366_ _0666_ clknet_leaf_65_clk_i memory\[14\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5578_ _2172_ _2179_ _2184_ _2189_ _1952_ _2190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_14_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3943__I1 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7134__I1 _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8297_ _0597_ clknet_leaf_128_clk_i net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4529_ _1475_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7317_ _3647_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6098__A1 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5623__C _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7248_ _1160_ memory\[8\]\[30\] _3577_ _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5145__I0 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6719__C _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_8_0_clk_i clknet_0_clk_i clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5845__B2 _2450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7611__S _3795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7179_ _3574_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_37_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7410__I _3685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6270__A1 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6022__B2 _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6470__B _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7058__S _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_46_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_136_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6897__S _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6325__A2 _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5136__I0 _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6089__A1 _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4210__S _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_170_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput9 data_i[12] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6137__S _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5041__S _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6261__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6364__C _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6013__A1 _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3900_ net6 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4880_ _1076_ memory\[25\]\[24\] _1660_ _1665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4880__S _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3870__I0 _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5775__I _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_95_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6550_ _2784_ memory\[0\]\[26\] _3141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_27_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5501_ memory\[22\]\[4\] _2114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_125_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6481_ _2848_ memory\[27\]\[25\] _3072_ _2850_ _3073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_112_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8220_ _0520_ clknet_leaf_12_clk_i memory\[28\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5432_ _2044_ _2046_ _1950_ _2047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8151_ _0451_ clknet_leaf_10_clk_i memory\[26\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5363_ memory\[12\]\[1\] memory\[13\]\[1\] _1978_ _1979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4314_ _1068_ memory\[17\]\[20\] _1358_ _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7102_ memory\[31\]\[25\] _1223_ _3528_ _3534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5827__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8082_ _0382_ clknet_leaf_43_clk_i memory\[24\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5294_ _1910_ _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4245_ _1299_ _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7033_ memory\[13\]\[25\] _1223_ _3491_ _3497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4176_ _1072_ memory\[15\]\[22\] _1280_ _1283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6252__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7935_ _0235_ clknet_leaf_172_clk_i memory\[1\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6004__A1 _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3861__I0 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7866_ _0166_ clknet_leaf_188_clk_i memory\[17\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6817_ _3382_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_102_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5685__I _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6555__A2 _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7797_ _0097_ clknet_leaf_195_clk_i memory\[15\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6748_ _1873_ _3333_ _2961_ _3334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6679_ _2884_ _3266_ _1913_ _3267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_131_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6510__S _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8418_ _0718_ clknet_leaf_156_clk_i memory\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5634__B _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8349_ _0649_ clknet_leaf_169_clk_i memory\[9\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5126__S _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5818__A1 _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6491__B2 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6465__B _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7291__I0 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6243__A1 _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_117_clk_i_I clknet_4_14_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5528__C _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4004__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7516__S _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4939__I _1673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5109__I0 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__I1 _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5809__A1 _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6482__A1 _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5285__A2 _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4030_ _1184_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6234__A1 _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5981_ _2208_ memory\[18\]\[14\] _2584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_59_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4932_ _1692_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7720_ _0020_ clknet_leaf_124_clk_i memory\[19\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_72_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7651_ memory\[6\]\[27\] net25 _3817_ _3825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4863_ _1273_ memory\[25\]\[16\] _1649_ _1656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4548__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4115__S _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7585__I1 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6602_ _3176_ _3181_ _3186_ _3191_ _2894_ _3192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_28_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4794_ _1619_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7582_ _3788_ _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6533_ memory\[23\]\[26\] _2713_ _3123_ _2006_ _3124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6464_ _2779_ _3056_ _2643_ _3057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8203_ _0503_ clknet_leaf_73_clk_i memory\[28\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5454__B _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5415_ _1909_ _2028_ _2029_ _2030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6395_ memory\[24\]\[23\] _2799_ _2989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5346_ _1877_ memory\[28\]\[1\] _1962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_11_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8134_ _0434_ clknet_leaf_163_clk_i memory\[26\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4785__S _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8065_ _0365_ clknet_leaf_175_clk_i memory\[24\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5277_ _1893_ _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4228_ _1313_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7016_ memory\[13\]\[17\] _1206_ _3480_ _3488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5276__A2 _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6473__A1 _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input28_I data_i[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4159_ _1272_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_104_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7918_ _0218_ clknet_leaf_99_clk_i memory\[1\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6505__S _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7849_ _0149_ clknet_leaf_87_clk_i memory\[17\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7336__S _3650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3864__S _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6179__C _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_43_clk_i_I clknet_4_4_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6839__I0 _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7071__S _3517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6464__A1 _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7264__I0 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6216__B2 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6519__A2 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6214__I _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 data_i[15] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_126_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4250__I0 _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput34 data_i[6] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7246__S _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput23 data_i[25] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_77_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5274__B _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5200_ _1127_ memory\[30\]\[14\] _1830_ _1835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_110_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6180_ _1872_ _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4553__I1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5131_ _1798_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5062_ _1267_ memory\[28\]\[13\] _1758_ _1762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4013_ net17 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_35_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6207__A1 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3949__S _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8752_ _1052_ clknet_leaf_70_clk_i memory\[7\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5964_ _2330_ net43 _2568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7703_ _0003_ clknet_leaf_192_clk_i memory\[7\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5895_ memory\[12\]\[12\] memory\[13\]\[12\] _2453_ _2500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7558__I1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8683_ _0983_ clknet_leaf_91_clk_i memory\[5\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4915_ _1683_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_23_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7634_ memory\[6\]\[19\] net16 _3806_ _3816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_62_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4846_ _1256_ memory\[25\]\[8\] _1638_ _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7565_ _3779_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4241__I0 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4777_ _1610_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6516_ _2938_ _2939_ memory\[5\]\[25\] _3108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_132_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7496_ _3742_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6447_ memory\[22\]\[24\] _3040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6995__S _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4544__I1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6694__A1 _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6378_ _2970_ _2972_ _2880_ _2973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8117_ _0417_ clknet_leaf_14_clk_i memory\[25\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5329_ _1930_ memory\[6\]\[0\] _1946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5404__S _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8048_ _0348_ clknet_leaf_51_clk_i memory\[23\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7246__I0 _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6462__C _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5421__A2 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5359__B _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7066__S _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4783__I1 _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6685__A1 _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7485__I0 _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4299__I0 _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4471__I0 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5680_ memory\[30\]\[8\] memory\[31\]\[8\] _2066_ _2289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_84_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4700_ _1250_ memory\[23\]\[5\] _1562_ _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_84_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4631_ _1530_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7350_ _3665_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4562_ _1493_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4774__I1 _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7281_ _1125_ memory\[3\]\[13\] _3625_ _3629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6301_ memory\[24\]\[21\] _2799_ _2897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4493_ _1456_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_122_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4526__I1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6232_ _2776_ memory\[11\]\[19\] _2829_ _2640_ _2830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_12_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6676__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6163_ memory\[23\]\[18\] _2713_ _2761_ _2671_ _2762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6094_ memory\[4\]\[16\] _2468_ _2695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7476__I0 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5114_ _1789_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5451__C _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5045_ _1250_ memory\[28\]\[5\] _1747_ _1753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7228__I0 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5651__A2 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__I _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6996_ _3477_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5947_ _2362_ memory\[10\]\[13\] _2551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8735_ _1035_ clknet_leaf_179_clk_i memory\[6\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6600__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8666_ _0966_ clknet_leaf_213_clk_i memory\[10\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5907__B _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5878_ _2108_ memory\[28\]\[12\] _2483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7617_ _3807_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7400__I0 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5693__I _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4214__I0 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4829_ _1637_ _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_63_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8597_ _0897_ clknet_leaf_187_clk_i memory\[4\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4303__S _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7548_ memory\[5\]\[10\] net7 _3770_ _3771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7479_ _1118_ memory\[10\]\[10\] _3733_ _3734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_216_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4517__I1 _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4102__I net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5134__S _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6419__A1 _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4973__S _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output59_I net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7219__I0 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_123_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__C _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3851__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5330__A1 _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7458__I0 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4692__I0 _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6383__B _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6850_ _3400_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5801_ memory\[15\]\[10\] _2357_ _2407_ _2307_ _2408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_76_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6781_ _1102_ memory\[9\]\[2\] _3361_ _3364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4444__I0 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8520_ _0820_ clknet_leaf_115_clk_i memory\[8\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5732_ _2108_ memory\[28\]\[9\] _2340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_58_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3993_ _1157_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_165_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5663_ _2269_ _2272_ _1950_ _2273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8451_ _0751_ clknet_leaf_136_clk_i memory\[31\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5219__S _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7402_ _1110_ memory\[0\]\[6\] _3686_ _3693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4614_ _1520_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8382_ _0682_ clknet_leaf_197_clk_i memory\[14\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5594_ _1879_ _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7333_ _3656_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4545_ _1483_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6649__A1 _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7434__S _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7264_ _1108_ memory\[3\]\[5\] _3614_ _3620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4476_ _1446_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6215_ memory\[20\]\[19\] memory\[21\]\[19\] _2812_ _2813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7195_ _3583_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5321__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6146_ _2330_ net47 _2746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5889__S _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4793__S _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6077_ _2629_ _2677_ _2495_ _2678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input10_I data_i[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ _1743_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4592__I _1486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_4_0_clk_i clknet_0_clk_i clknet_4_4_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5388__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7609__S _3795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6979_ _1167_ _1485_ _3468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_200_clk_i clknet_4_2_0_clk_i clknet_leaf_200_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8718_ _1018_ clknet_leaf_68_clk_i memory\[6\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8649_ _0949_ clknet_leaf_112_clk_i memory\[10\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3936__I _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5356__C _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_6_clk_i clknet_4_1_0_clk_i clknet_leaf_6_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_11_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_215_clk_i clknet_4_0_0_clk_i clknet_leaf_215_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7688__I0 _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_56_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5863__A2 _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6187__C _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4208__S _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5379__A1 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5918__A3 _2521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4977__I1 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5039__S _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4878__S _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7254__S _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4330_ _1084_ memory\[17\]\[28\] _1358_ _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6378__B _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4261_ _1330_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6000_ _2418_ _2601_ _2602_ _2603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_91_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I address_i[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4192_ _1089_ memory\[15\]\[30\] _1239_ _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5502__S _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5606__A2 _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7951_ _0251_ clknet_leaf_51_clk_i memory\[20\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7882_ _0182_ clknet_leaf_86_clk_i memory\[18\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5301__I _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4118__S _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6902_ _3427_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6833_ _1154_ memory\[9\]\[27\] _3383_ _3391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7429__S _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4417__I0 _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6560__C _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6764_ _3347_ _3349_ _1916_ _3350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3976_ net21 _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_134_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5715_ memory\[4\]\[8\] _1998_ _2324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6695_ _2000_ memory\[29\]\[30\] _3281_ _1925_ _3282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8503_ _0803_ clknet_leaf_209_clk_i memory\[11\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_98_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8434_ _0734_ clknet_leaf_75_clk_i memory\[13\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5646_ _2253_ _2255_ _1916_ _2256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_116_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8365_ _0665_ clknet_leaf_65_clk_i memory\[14\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5577_ _1997_ _2185_ _2187_ _2188_ _2189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5971__I _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5542__A1 _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7164__S _3564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4528_ memory\[20\]\[22\] _1217_ _1472_ _1475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8296_ _0596_ clknet_leaf_120_clk_i net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7316_ _1160_ memory\[3\]\[30\] _3613_ _3647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7247_ _3610_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4459_ _1072_ memory\[1\]\[22\] _1435_ _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6893__I1 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3856__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7047__A1 _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7178_ memory\[11\]\[29\] _1231_ _3564_ _3574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6129_ _2310_ memory\[11\]\[17\] _2728_ _2640_ _2729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_99_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A2 _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4408__I0 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3867__S _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5081__I0 _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5781__A1 _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7138__I _3541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_154_clk_i clknet_4_10_0_clk_i clknet_leaf_154_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5533__A1 _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4698__S _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_169_clk_i clknet_4_8_0_clk_i clknet_leaf_169_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_31_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_113_clk_i_I clknet_4_14_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6884__I1 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_107_clk_i clknet_4_15_0_clk_i clknet_leaf_107_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_82_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6013__A2 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5072__I0 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_38_clk_i_I clknet_4_4_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5772__A1 _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5500_ _2110_ _2112_ _1890_ _2113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6480_ _2898_ memory\[26\]\[25\] _3072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5524__A1 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5431_ _1941_ _2045_ _1994_ _2046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8150_ _0450_ clknet_leaf_11_clk_i memory\[26\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5362_ _1884_ _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8081_ _0381_ clknet_leaf_49_clk_i memory\[24\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4313_ _1335_ _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7101_ _3533_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5293_ _1059_ _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_10_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7032_ _3496_ _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4244_ _1321_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4886__I0 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4175_ _1282_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_3_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7934_ _0234_ clknet_leaf_171_clk_i memory\[1\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7865_ _0165_ clknet_leaf_20_clk_i memory\[17\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6571__B _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_71_clk_i clknet_4_7_0_clk_i clknet_leaf_71_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6816_ _1137_ memory\[9\]\[19\] _3372_ _3382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7796_ _0096_ clknet_leaf_28_clk_i memory\[15\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7052__I1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5763__A1 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6747_ memory\[16\]\[31\] memory\[17\]\[31\] _1885_ _3333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3959_ _1134_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6678_ memory\[2\]\[29\] memory\[3\]\[29\] _1911_ _3266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_21_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6797__I _3360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_86_clk_i clknet_4_12_0_clk_i clknet_leaf_86_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5515__A1 _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8417_ _0717_ clknet_leaf_151_clk_i memory\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5629_ _1871_ _2060_ memory\[25\]\[7\] _2239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_103_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4311__S _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8348_ _0648_ clknet_leaf_206_clk_i memory\[9\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_131_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7622__S _3806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8279_ _0579_ clknet_leaf_18_clk_i memory\[30\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6866__I1 _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5142__S _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6238__S _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6491__A2 _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_24_clk_i clknet_4_3_0_clk_i clknet_leaf_24_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4981__S _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4006__A1 _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_39_clk_i clknet_4_4_0_clk_i clknet_leaf_39_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_64_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_1_Left_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7043__I1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5506__A1 _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6656__B _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6857__I1 _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6482__A2 _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6375__C _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5980_ _2580_ _2294_ _2582_ _2250_ _2583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_63_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4931_ _1273_ memory\[26\]\[16\] _1685_ _1692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4862_ _1655_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7650_ _3824_ _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5045__I0 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6601_ _2933_ _3187_ _3189_ _3190_ _3191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4793_ memory\[24\]\[15\] _1202_ _1613_ _1619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6793__I0 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5745__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7581_ memory\[5\]\[26\] net24 _3781_ _3788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6532_ memory\[20\]\[26\] memory\[21\]\[26\] _2812_ _3123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5735__B _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ memory\[8\]\[24\] memory\[9\]\[24\] _2780_ _3056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8202_ _0502_ clknet_leaf_131_clk_i memory\[28\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5414_ _1057_ _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5227__S _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4020__I1 _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8133_ _0433_ clknet_leaf_164_clk_i memory\[26\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6394_ _2846_ _2964_ _2987_ _2988_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__7442__S _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5345_ _1857_ _1956_ _1959_ _1960_ _1961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__4859__I0 _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5276_ _1295_ _1060_ _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_8064_ _0364_ clknet_leaf_133_clk_i memory\[23\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7015_ _3487_ _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4227_ _1263_ memory\[29\]\[11\] _1311_ _1313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4158_ _1271_ memory\[15\]\[15\] _1261_ _1272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ _1224_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7917_ _0217_ clknet_leaf_99_clk_i memory\[1\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5984__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7025__I1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7848_ _0148_ clknet_leaf_125_clk_i memory\[17\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7779_ _0079_ clknet_leaf_156_clk_i memory\[15\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4105__I net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5645__B _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_115_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4011__I1 _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5380__B _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5600__S _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6216__A2 _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7016__I1 _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4216__S _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7527__S _3759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5727__A1 _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 data_i[16] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_115_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput35 data_i[7] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5555__B _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput24 data_i[26] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5047__S _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3854__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6230__I _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6152__A1 _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7262__S _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4886__S _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5130_ _1267_ memory\[2\]\[13\] _1794_ _1798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5061_ _1761_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4012_ _1172_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4069__I1 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5963_ _2550_ _2555_ _2560_ _2566_ _2428_ _2567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_8751_ _1051_ clknet_leaf_68_clk_i memory\[7\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_88_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4914_ _1256_ memory\[26\]\[8\] _1674_ _1683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7702_ _0002_ clknet_leaf_188_clk_i memory\[7\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5894_ memory\[14\]\[12\] _2499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_118_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8682_ _0982_ clknet_leaf_85_clk_i memory\[5\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5718__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7633_ _3815_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4845_ _1646_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7564_ memory\[5\]\[18\] net15 _3770_ _3779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4776_ memory\[24\]\[7\] _1185_ _1602_ _1610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6391__A1 _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5465__B _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6515_ _2981_ memory\[7\]\[25\] _3106_ _2983_ _3107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_114_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7495_ _1135_ memory\[10\]\[18\] _3733_ _3742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6143__A1 _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6446_ _3036_ _3038_ _2757_ _3039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7172__S _3564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6377_ _2779_ _2971_ _2643_ _2972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8116_ _0416_ clknet_leaf_35_clk_i memory\[25\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5328_ _1857_ _1942_ _1943_ _1944_ _1945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA_clkbuf_leaf_7_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8047_ _0347_ clknet_leaf_51_clk_i memory\[23\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5259_ _1861_ _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_3_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_212_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3939__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7347__S _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_91_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6134__A1 _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5822__C _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6437__A2 _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6426__S _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6653__C _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5948__A1 _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6225__I _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4630_ memory\[22\]\[5\] _1181_ _1524_ _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4561_ memory\[21\]\[5\] _1181_ _1487_ _1493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6300_ _2846_ _2870_ _2895_ _2896_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7280_ _3628_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4492_ memory\[20\]\[5\] _1181_ _1450_ _1456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6231_ _2828_ memory\[10\]\[19\] _2829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_110_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6162_ memory\[20\]\[18\] memory\[21\]\[18\] _2346_ _2761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_161_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5113_ _1250_ memory\[2\]\[5\] _1783_ _1789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6093_ _2691_ _2693_ _2421_ _2694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_85_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5304__I _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5044_ _1752_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6995_ memory\[13\]\[7\] _1185_ _3469_ _3477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_137_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ _2547_ _2406_ _2549_ _2360_ _2550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_47_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8734_ _1034_ clknet_leaf_196_clk_i memory\[6\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6600__A2 _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5877_ _2332_ _2478_ _2480_ _2481_ _2482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_48_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8665_ _0965_ clknet_leaf_212_clk_i memory\[10\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7616_ memory\[6\]\[10\] net7 _3806_ _3807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_86_clk_i_I clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4828_ _1298_ _1599_ _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_62_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8596_ _0896_ clknet_leaf_80_clk_i memory\[4\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6364__A1 _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7547_ _3758_ _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4759_ _1598_ _1599_ _1600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7478_ _3721_ _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_8_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6429_ memory\[4\]\[23\] _2934_ _3023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_0_0_clk_i clknet_0_clk_i clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_128_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7630__S _3806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6473__C _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7077__S _3517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6355__A1 _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6107__A1 _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6156__S _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6664__B _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5060__S _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6969__I0 _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_108_clk_i_I clknet_4_15_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7630__I1 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5800_ memory\[12\]\[10\] memory\[13\]\[10\] _1978_ _2407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6780_ _3363_ _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3992_ memory\[19\]\[28\] _1156_ _1140_ _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5397__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5731_ _2332_ _2334_ _2336_ _2338_ _2339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_73_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4404__S _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5662_ _1941_ _2271_ _2136_ _2272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8450_ _0750_ clknet_leaf_135_clk_i memory\[31\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7394__I0 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6346__A1 _2922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7401_ _3692_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4613_ memory\[21\]\[30\] _1233_ _1486_ _1520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8381_ _0681_ clknet_leaf_197_clk_i memory\[14\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5593_ memory\[20\]\[6\] memory\[21\]\[6\] _1897_ _2204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_130_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7332_ _1108_ memory\[4\]\[5\] _3650_ _3656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4544_ memory\[20\]\[30\] _1233_ _1449_ _1483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4203__I _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7263_ _3619_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_96_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6214_ _1059_ _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4475_ _1089_ memory\[1\]\[30\] _1412_ _1446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5235__S _1818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7194_ _1106_ memory\[8\]\[4\] _3578_ _3583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5462__C _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5872__A3 _2476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6145_ _2727_ _2732_ _2739_ _2744_ _2428_ _2745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_96_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5034__I _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7450__S _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6076_ memory\[16\]\[16\] memory\[17\]\[16\] _2630_ _2677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5027_ memory\[27\]\[29\] _1231_ _1733_ _1743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8717_ _1017_ clknet_leaf_91_clk_i memory\[6\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6978_ _3467_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6585__B2 _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5929_ memory\[30\]\[13\] memory\[31\]\[13\] _2532_ _2533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8648_ _0948_ clknet_leaf_115_clk_i memory\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4314__S _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8579_ _0879_ clknet_leaf_120_clk_i memory\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6749__B _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5560__A2 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5145__S _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4371__I0 _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4674__I1 _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5547__C _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6328__A1 _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7376__I0 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7535__S _3759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4260_ _1082_ memory\[29\]\[27\] _1322_ _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4362__I0 _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_34_clk_i_I clknet_4_4_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4894__S _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4191_ _1290_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7270__S _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7300__I0 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7950_ _0250_ clknet_leaf_52_clk_i memory\[20\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7881_ _0181_ clknet_leaf_127_clk_i memory\[18\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6901_ memory\[14\]\[27\] _1227_ _3419_ _3427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6832_ _3390_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_18_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6567__A1 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3975_ _1145_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6763_ _1883_ _3348_ _1913_ _3349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_128_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5790__A2 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5714_ _2320_ _2322_ _1950_ _2323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6694_ _2001_ memory\[28\]\[30\] _3281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6319__A1 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8502_ _0802_ clknet_leaf_208_clk_i memory\[11\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8433_ _0733_ clknet_leaf_58_clk_i memory\[13\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5645_ _2163_ _2254_ _2029_ _2255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_98_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8364_ _0664_ clknet_leaf_65_clk_i memory\[14\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5576_ _2005_ _2007_ memory\[5\]\[5\] _2188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_60_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8295_ _0595_ clknet_leaf_123_clk_i net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4527_ _1474_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7315_ _3646_ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7246_ _1158_ memory\[8\]\[29\] _3600_ _3610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4458_ _1437_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7177_ _3573_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6128_ _2362_ memory\[10\]\[17\] _2728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4389_ _1400_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3856__A2 _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7180__S _3541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6059_ _2382_ memory\[27\]\[16\] _2659_ _2384_ _2660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_99_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4309__S _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6558__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6323__I _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5367__C _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4979__S _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7355__S _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6730__A1 _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5297__A1 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4344__I0 _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_69_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4647__I1 _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3857__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7349__I0 _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5430_ memory\[2\]\[2\] memory\[3\]\[2\] _1992_ _2045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6721__A1 _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_10_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5361_ memory\[14\]\[1\] _1977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8080_ _0380_ clknet_leaf_49_clk_i memory\[24\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_93_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4312_ _1357_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5292_ _1872_ _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7100_ memory\[31\]\[24\] _1221_ _3528_ _3533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4243_ _1056_ memory\[29\]\[19\] _1311_ _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7031_ memory\[13\]\[24\] _1221_ _3491_ _3496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4174_ _1070_ memory\[15\]\[21\] _1280_ _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5312__I _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_5_clk_i clknet_4_1_0_clk_i clknet_leaf_5_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4638__I1 _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_214_clk_i clknet_4_0_0_clk_i clknet_leaf_214_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7933_ _0233_ clknet_leaf_196_clk_i memory\[1\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5460__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3968__S _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7864_ _0164_ clknet_leaf_21_clk_i memory\[17\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6815_ _3381_ _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7795_ _0095_ clknet_leaf_79_clk_i memory\[15\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_4_7_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6746_ _1876_ memory\[19\]\[31\] _3331_ _2003_ _3332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_19_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3958_ memory\[19\]\[17\] _1133_ _1119_ _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4799__S _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4810__I1 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6677_ _1904_ memory\[1\]\[29\] _3264_ _2975_ _3265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3889_ _1085_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8416_ _0716_ clknet_leaf_181_clk_i memory\[16\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5628_ _1862_ memory\[27\]\[7\] _2237_ _1867_ _2238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_5_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8347_ _0647_ clknet_leaf_214_clk_i memory\[9\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5559_ memory\[15\]\[5\] _1922_ _2170_ _1925_ _2171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_131_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5931__B _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8278_ _0578_ clknet_leaf_19_clk_i memory\[30\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4326__I0 _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7512__I0 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6746__C _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7229_ _3601_ _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_69_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5451__A1 _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6481__C _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4801__I1 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7085__S _3517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6703__A1 _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_207_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5560__C _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5690__A1 _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6228__I _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5442__A1 _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4930_ _1691_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_111_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4861_ _1271_ memory\[25\]\[15\] _1649_ _1655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6600_ _2938_ _2939_ memory\[5\]\[27\] _3190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4792_ _1618_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7580_ _3787_ _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6531_ memory\[22\]\[26\] _3122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6462_ _2776_ memory\[11\]\[24\] _3054_ _2640_ _3055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_112_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8201_ _0501_ clknet_leaf_127_clk_i memory\[28\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5413_ memory\[16\]\[2\] memory\[17\]\[2\] _1911_ _2028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6393_ _2796_ net53 _2988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_120_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8132_ _0432_ clknet_leaf_164_clk_i memory\[26\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5344_ _1871_ _1873_ memory\[25\]\[1\] _1960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_112_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8063_ _0363_ clknet_leaf_132_clk_i memory\[23\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5275_ memory\[22\]\[0\] _1892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7014_ memory\[13\]\[16\] _1204_ _3480_ _3487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4226_ _1312_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5470__C _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4157_ net12 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5681__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_153_clk_i clknet_4_10_0_clk_i clknet_leaf_153_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_128_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4088_ memory\[12\]\[25\] _1223_ _1213_ _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7916_ _0216_ clknet_leaf_105_clk_i memory\[1\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_104_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7847_ _0147_ clknet_leaf_124_clk_i memory\[17\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_168_clk_i clknet_4_8_0_clk_i clknet_leaf_168_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_3_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6802__S _3372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_156_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7778_ _0078_ clknet_leaf_156_clk_i memory\[15\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6729_ _1854_ net62 _3316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4322__S _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3960__I net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__S _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6476__C _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4992__S _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5027__I1 _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput14 data_i[17] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput36 data_i[8] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput25 data_i[27] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_134_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7543__S _3759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4031__I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5360__B1 _1970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5571__B _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7342__I _3649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4966__I _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_70_clk_i clknet_4_7_0_clk_i clknet_leaf_70_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5060_ _1265_ memory\[28\]\[12\] _1758_ _1761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5998__S _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4011_ memory\[12\]\[0\] _1164_ _1171_ _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5415__A1 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5962_ _2467_ _2561_ _2564_ _2565_ _2566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_8750_ _1050_ clknet_leaf_68_clk_i memory\[7\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_85_clk_i clknet_4_12_0_clk_i clknet_leaf_85_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5966__A2 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4913_ _1682_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7701_ _0001_ clknet_leaf_187_clk_i memory\[7\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5893_ _2482_ _2487_ _2491_ _2497_ _2403_ _2498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_8681_ _0981_ clknet_leaf_110_clk_i memory\[5\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5718__A2 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7632_ memory\[6\]\[18\] net15 _3806_ _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4844_ _1254_ memory\[25\]\[7\] _1638_ _1646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5746__B _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7563_ _3778_ _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4775_ _1609_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6514_ _1864_ memory\[6\]\[25\] _3106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7494_ _3741_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_23_clk_i clknet_4_6_0_clk_i clknet_leaf_23_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6143__A2 _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6445_ _2754_ _3037_ _2666_ _3038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6376_ memory\[8\]\[22\] memory\[9\]\[22\] _2780_ _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6069__S _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8115_ _0415_ clknet_leaf_44_clk_i memory\[25\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5327_ memory\[3\]\[0\] _1922_ _1858_ memory\[0\]\[0\] _1944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8046_ _0346_ clknet_leaf_52_clk_i memory\[23\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_82_clk_i_I clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_38_clk_i clknet_4_4_0_clk_i clknet_leaf_38_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input33_I data_i[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5258_ _1857_ _1860_ _1868_ _1874_ _1875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5189_ _1116_ memory\[30\]\[9\] _1819_ _1829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4209_ _1303_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_3_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__A2 _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7628__S _3806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5009__I1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6532__S _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5656__B _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5375__C _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7182__I1 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6487__B _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5893__B2 _2497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4940__I0 _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5645__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4227__S _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5566__B _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5058__S _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4560_ _1492_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5285__C _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6373__A2 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4491_ _1455_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6230_ _1869_ _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_leaf_104_clk_i_I clknet_4_15_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4931__I0 _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6161_ _1893_ _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5112_ _1788_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6092_ _2418_ _2692_ _2602_ _2693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5043_ _1248_ memory\[28\]\[4\] _1747_ _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_0_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6061__A1 _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5320__I _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6987__I1 _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6994_ _3476_ _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5945_ memory\[15\]\[13\] _2357_ _2548_ _2307_ _2549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_125_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7448__S _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8733_ _1033_ clknet_leaf_195_clk_i memory\[6\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5876_ _2337_ _2060_ memory\[25\]\[12\] _2481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_91_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_29_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8664_ _0964_ clknet_leaf_211_clk_i memory\[10\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7615_ _3794_ _3806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4827_ _1636_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8595_ _0895_ clknet_leaf_83_clk_i memory\[4\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7546_ _3769_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4758_ net3 _1165_ _1094_ _1599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_44_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7477_ _3732_ _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4689_ _1561_ _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_44_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7164__I1 _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5175__I0 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6428_ _3019_ _3021_ _2887_ _3022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5875__A1 _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6359_ memory\[22\]\[22\] _2954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5627__A1 _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8029_ _0329_ clknet_leaf_36_clk_i memory\[22\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6754__C _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6052__A1 _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7155__I1 _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3964__I1 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6680__B _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3991_ net26 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_29_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7268__S _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_30_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5730_ _2337_ _2060_ memory\[25\]\[9\] _2338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_33_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5661_ memory\[2\]\[7\] memory\[3\]\[7\] _2270_ _2271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7400_ _1108_ memory\[0\]\[5\] _3686_ _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4612_ _1519_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8380_ _0680_ clknet_leaf_0_clk_i memory\[14\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5592_ memory\[22\]\[6\] _2203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3955__I1 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7331_ _3655_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4543_ _1482_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5743__C _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7262_ _1106_ memory\[3\]\[4\] _3614_ _3619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5157__I0 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5857__A1 _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6213_ memory\[22\]\[19\] _2811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4904__I0 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4474_ _1445_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7193_ _3582_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5315__I _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5609__A1 _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6144_ _2467_ _2740_ _2742_ _2743_ _2744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6075_ _2626_ memory\[19\]\[16\] _2675_ _2541_ _2676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5026_ _1742_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6282__A1 _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6977_ _1162_ memory\[16\]\[31\] _3432_ _3467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6590__B _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8716_ _1016_ clknet_leaf_90_clk_i memory\[6\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5928_ _1884_ _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_76_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7178__S _3564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6585__A2 _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5859_ _2418_ _2464_ _2136_ _2465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8647_ _0947_ clknet_leaf_115_clk_i memory\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6810__S _3372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8578_ _0878_ clknet_leaf_120_clk_i memory\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3946__I1 _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7529_ memory\[5\]\[1\] net17 _3759_ _3761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5653__C _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4330__S _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7641__S _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5161__S _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6025__A1 _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3882__I0 _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4505__S _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6576__A2 _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5828__C _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4339__A1 _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6720__S _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5844__B _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3937__I1 _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5563__C _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7128__I1 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7615__I _3794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6675__B _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4190_ _1086_ memory\[15\]\[29\] _1280_ _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6167__S _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7880_ _0180_ clknet_leaf_125_clk_i memory\[18\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6900_ _3426_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3873__I0 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6016__A1 _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6831_ _1152_ memory\[9\]\[26\] _3383_ _3390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_18_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4415__S _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3974_ memory\[19\]\[22\] _1144_ _1140_ _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8501_ _0801_ clknet_leaf_198_clk_i memory\[11\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6762_ memory\[2\]\[31\] memory\[3\]\[31\] _1911_ _3348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5713_ _1941_ _2321_ _2136_ _2322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6693_ _1887_ _3276_ _3278_ _3279_ _3280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_57_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8432_ _0732_ clknet_leaf_60_clk_i memory\[13\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5644_ memory\[16\]\[7\] memory\[17\]\[7\] _2164_ _2254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_98_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8363_ _0663_ clknet_leaf_77_clk_i memory\[14\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5575_ _2049_ memory\[7\]\[5\] _2186_ _2051_ _2187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6569__C _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7314_ _1158_ memory\[3\]\[29\] _3636_ _3646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4526_ memory\[20\]\[21\] _1215_ _1472_ _1474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8294_ _0594_ clknet_leaf_120_clk_i net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_133_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7245_ _3609_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4457_ _1070_ memory\[1\]\[21\] _1435_ _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7176_ memory\[11\]\[28\] _1229_ _3564_ _3573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6127_ _2724_ _2406_ _2726_ _2360_ _2727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4388_ _1070_ memory\[18\]\[21\] _1398_ _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6255__A1 _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6058_ _2432_ memory\[26\]\[16\] _2659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_134_Right_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5009_ memory\[27\]\[20\] _1212_ _1733_ _1734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3864__I0 _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6802__I0 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6558__A2 _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4060__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3963__I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_15_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6494__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6715__S _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_203_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4235__S _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4280__I0 _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4034__I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5066__S _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6721__A2 _3307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6389__C _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_33_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5360_ _1961_ _1966_ _1970_ _1975_ _1918_ _1976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_112_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4311_ _1056_ memory\[17\]\[19\] _1347_ _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5291_ _1904_ memory\[19\]\[0\] _1906_ _1907_ _1908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7281__S _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4242_ _1320_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_4_14_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6485__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7030_ _3495_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6237__A1 _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4173_ _1281_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7285__I0 _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_42_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7932_ _0232_ clknet_leaf_197_clk_i memory\[1\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7863_ _0163_ clknet_leaf_23_clk_i memory\[17\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7794_ _0094_ clknet_leaf_75_clk_i memory\[15\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ _1135_ memory\[9\]\[18\] _3372_ _3381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3957_ net14 _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_92_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6745_ _1877_ memory\[18\]\[31\] _3331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_102_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6360__S _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8415_ _0715_ clknet_leaf_182_clk_i memory\[16\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6676_ _1905_ memory\[0\]\[29\] _3264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3888_ _1084_ memory\[7\]\[28\] _1066_ _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5627_ _1957_ memory\[26\]\[7\] _2237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6712__A2 _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4574__I1 _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8346_ _0646_ clknet_leaf_213_clk_i memory\[9\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5558_ memory\[12\]\[5\] memory\[13\]\[5\] _1978_ _2170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4509_ memory\[20\]\[13\] _1198_ _1461_ _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8277_ _0577_ clknet_leaf_189_clk_i memory\[30\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5489_ _1855_ _2080_ _2101_ _2102_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_53_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7228_ _1139_ memory\[8\]\[20\] _3600_ _3601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_152_clk_i_I clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7159_ _3541_ _3564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_69_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7579__I1 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6400__A1 _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_77_clk_i_I clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4262__I0 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7366__S _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7200__I0 _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4565__I1 _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6467__A1 _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5841__C _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6219__A1 _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6672__C _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4860_ _1654_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_28_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4791_ memory\[24\]\[14\] _1200_ _1613_ _1618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6530_ _3118_ _3120_ _2757_ _3121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6461_ _2828_ memory\[10\]\[24\] _3054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8200_ _0500_ clknet_leaf_128_clk_i memory\[28\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5412_ _1904_ memory\[19\]\[2\] _2026_ _1907_ _2027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6392_ _2968_ _2973_ _2979_ _2986_ _2894_ _2987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_30_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8131_ _0431_ clknet_leaf_165_clk_i memory\[26\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5343_ _1862_ memory\[27\]\[1\] _1958_ _1867_ _1959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_63_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8062_ _0362_ clknet_leaf_23_clk_i memory\[23\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5274_ _1881_ _1888_ _1890_ _1891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7013_ _3486_ _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4225_ _1260_ memory\[29\]\[10\] _1311_ _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4156_ _1270_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7258__I0 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5433__A2 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6582__C _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6630__A1 _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4087_ net23 _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7915_ _0215_ clknet_leaf_103_clk_i memory\[1\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_104_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5479__B _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7846_ _0146_ clknet_leaf_126_clk_i memory\[17\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4989_ _1723_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7186__S _3578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7777_ _0077_ clknet_leaf_151_clk_i memory\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4795__I1 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4603__S _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6728_ _3299_ _3304_ _3309_ _3314_ _1063_ _3315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6659_ memory\[23\]\[29\] _1895_ _3246_ _2006_ _3247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_33_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6697__A1 _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8329_ _0629_ clknet_leaf_88_clk_i memory\[9\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7497__I0 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6449__B2 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5672__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6492__C _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7421__I0 _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4235__I0 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7096__S _3528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4513__S _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput37 data_i[9] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput15 data_i[18] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_80_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput26 data_i[28] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_123_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4538__I1 _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_4_clk_i clknet_4_1_0_clk_i clknet_leaf_4_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_40_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_213_clk_i clknet_4_0_0_clk_i clknet_leaf_213_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4010_ _1170_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5961_ _2472_ _2473_ memory\[5\]\[13\] _2565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_88_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_100_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8680_ _0980_ clknet_leaf_110_clk_i memory\[5\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7700_ _0000_ clknet_leaf_27_clk_i memory\[7\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4912_ _1254_ memory\[26\]\[7\] _1674_ _1682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6903__S _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5892_ _2493_ _2496_ _2302_ _2497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7631_ _3814_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4843_ _1645_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7562_ memory\[5\]\[17\] net14 _3770_ _3778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4423__S _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4774_ memory\[24\]\[6\] _1183_ _1602_ _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7493_ _1133_ memory\[10\]\[17\] _3733_ _3741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6513_ memory\[4\]\[25\] _2934_ _3105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5318__I _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6444_ memory\[30\]\[24\] memory\[31\]\[24\] _1923_ _3037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6679__A1 _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6375_ _2776_ memory\[11\]\[22\] _2969_ _2640_ _2970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7479__I0 _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8114_ _0414_ clknet_leaf_43_clk_i memory\[25\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5326_ memory\[1\]\[0\] _1870_ _1909_ _1943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_11_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8045_ _0345_ clknet_leaf_53_clk_i memory\[23\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_25_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5257_ _1871_ _1873_ memory\[25\]\[0\] _1874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4208_ _1244_ memory\[29\]\[2\] _1300_ _1303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_110_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5188_ _1828_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input26_I data_i[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4139_ _1258_ memory\[15\]\[9\] _1240_ _1259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6603__A1 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4465__I0 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7829_ _0129_ clknet_leaf_22_clk_i memory\[29\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4768__I1 _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5590__A1 _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4132__I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5342__A1 _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4208__I0 _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4243__S _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7554__S _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_152_clk_i clknet_4_11_0_clk_i clknet_leaf_152_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_111_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4490_ memory\[20\]\[4\] _1179_ _1450_ _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_122_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5074__S _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3881__I net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6160_ memory\[22\]\[18\] _2759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6397__C _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5111_ _1248_ memory\[2\]\[4\] _1783_ _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_167_clk_i clknet_4_8_0_clk_i clknet_leaf_167_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6091_ memory\[2\]\[16\] memory\[3\]\[16\] _2270_ _2692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_199_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5042_ _1751_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6993_ memory\[13\]\[6\] _1183_ _3469_ _3476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5944_ memory\[12\]\[13\] memory\[13\]\[13\] _2453_ _2548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_105_clk_i clknet_4_15_0_clk_i clknet_leaf_105_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4998__I1 _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8732_ _1032_ clknet_leaf_3_clk_i memory\[6\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5875_ _2382_ memory\[27\]\[12\] _2479_ _2384_ _2480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_8_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8663_ _0963_ clknet_leaf_206_clk_i memory\[10\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8594_ _0894_ clknet_leaf_76_clk_i memory\[4\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7614_ _3805_ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4826_ memory\[24\]\[31\] _1235_ _1601_ _1636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7545_ memory\[5\]\[9\] net37 _3759_ _3769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4757_ _1597_ _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3992__S _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7464__S _3722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7476_ _1116_ memory\[10\]\[9\] _3722_ _3732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4688_ _1560_ _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_102_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6427_ _2884_ _3020_ _2602_ _3021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_112_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6358_ _2950_ _2952_ _2757_ _2953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_8_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ memory\[15\]\[0\] _1922_ _1924_ _1925_ _1926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6808__S _3372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5712__S _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6289_ _2884_ _2885_ _2602_ _2886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8028_ _0328_ clknet_leaf_37_clk_i memory\[22\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4328__S _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4438__I0 _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6052__A2 _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7639__S _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6770__C _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3966__I net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4063__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5159__S _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6342__I _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4998__S _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5563__A1 _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7374__S _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_84_clk_i clknet_4_12_0_clk_i clknet_leaf_84_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_99_clk_i clknet_4_13_0_clk_i clknet_leaf_99_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5618__A2 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6043__A2 _2644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4429__I0 _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4037__I net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_22_clk_i clknet_4_3_0_clk_i clknet_leaf_22_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6453__S _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3990_ _1155_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5660_ _1910_ _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_37_clk_i clknet_4_4_0_clk_i clknet_leaf_37_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4611_ memory\[21\]\[29\] _1231_ _1509_ _1519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5554__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5591_ _2198_ _2201_ _1890_ _2202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_13_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7330_ _1106_ memory\[4\]\[4\] _3650_ _3655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4542_ memory\[20\]\[29\] _1231_ _1472_ _1482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7261_ _3618_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4473_ _1086_ memory\[1\]\[29\] _1435_ _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_96_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6212_ _2807_ _2809_ _2757_ _2810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7192_ _1104_ memory\[8\]\[3\] _3578_ _3582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6143_ _2472_ _2473_ memory\[5\]\[17\] _2743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_127_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6074_ _2674_ memory\[18\]\[16\] _2675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5025_ memory\[27\]\[28\] _1229_ _1733_ _1742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6976_ _3466_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5093__I0 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5927_ _2529_ memory\[29\]\[13\] _2530_ _2389_ _2531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8715_ _1015_ clknet_leaf_84_clk_i memory\[6\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4840__I0 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5858_ memory\[2\]\[11\] memory\[3\]\[11\] _2270_ _2464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8646_ _0946_ clknet_leaf_116_clk_i memory\[10\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5789_ memory\[23\]\[10\] _2247_ _2395_ _2205_ _2396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7194__S _3578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8577_ _0877_ clknet_leaf_146_clk_i memory\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4809_ _1627_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4611__S _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7528_ _3760_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7459_ _3723_ _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6111__B _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_79_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3859__A1 _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5950__B _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6337__I _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output57_I net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7073__I1 _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_147_clk_i_I clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__A1 _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4521__S _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5839__A2 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_97_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4898__I0 _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6887__I1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5860__B _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6448__S _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5352__S _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7279__S _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7064__I1 _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6830_ _3389_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_18_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6761_ _1904_ memory\[1\]\[31\] _3346_ _2975_ _3347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5712_ memory\[2\]\[8\] memory\[3\]\[8\] _2270_ _2321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8500_ _0800_ clknet_leaf_27_clk_i memory\[11\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3973_ net20 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6692_ _1870_ _1990_ memory\[25\]\[30\] _3279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_127_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8431_ _0731_ clknet_leaf_62_clk_i memory\[13\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5643_ _2160_ memory\[19\]\[7\] _2252_ _2075_ _2253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5527__A1 _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5574_ _2096_ memory\[6\]\[5\] _2186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4431__S _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8362_ _0662_ clknet_leaf_178_clk_i memory\[14\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4525_ _1473_ _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7313_ _3645_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8293_ _0593_ clknet_leaf_120_clk_i net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_133_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6878__I1 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7244_ _1156_ memory\[8\]\[28\] _3600_ _3609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4456_ _1436_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4387_ _1399_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7175_ _3572_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6126_ memory\[15\]\[17\] _2357_ _2725_ _2307_ _2726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6255__A2 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6057_ memory\[24\]\[16\] _2333_ _2658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_107_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5008_ _1710_ _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_107_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5066__I0 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_120_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5766__A1 _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6959_ _1144_ memory\[16\]\[22\] _3455_ _3458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6821__S _3383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5518__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8629_ _0929_ clknet_leaf_197_clk_i memory\[0\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_73_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5900__S _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5839__C _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5855__B _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4032__I1 _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4050__I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7562__S _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4310_ _1356_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5290_ _1866_ _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4241_ _1277_ memory\[29\]\[18\] _1311_ _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5590__B _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4172_ _1068_ memory\[15\]\[20\] _1280_ _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5996__A1 _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7931_ _0231_ clknet_leaf_207_clk_i memory\[1\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7037__I1 _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7862_ _0162_ clknet_leaf_26_clk_i memory\[17\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6813_ _3380_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7793_ _0093_ clknet_leaf_70_clk_i memory\[15\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3956_ _1132_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6744_ _3327_ _1893_ _3329_ _1937_ _3330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_18_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6675_ _3260_ _3262_ _2880_ _3263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_135_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4161__S _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5484__C _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8414_ _0714_ clknet_leaf_186_clk_i memory\[16\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3887_ net26 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5626_ memory\[24\]\[7\] _1859_ _2236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4023__I1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5920__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7472__S _3722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8345_ _0645_ clknet_leaf_214_clk_i memory\[9\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5557_ memory\[14\]\[5\] _2169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4508_ _1464_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8276_ _0576_ clknet_leaf_31_clk_i memory\[30\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5488_ _1954_ net64 _2102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6596__B _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4439_ _1427_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7227_ _3577_ _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7158_ _3563_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6109_ memory\[30\]\[17\] memory\[31\]\[17\] _2532_ _2709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6816__S _3372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7089_ memory\[31\]\[19\] _1210_ _3517_ _3527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4336__S _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5659__C _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5039__I0 _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6787__I0 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7647__S _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4135__I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4411__A1 _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5167__S _1782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5394__C _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4014__I1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5911__A1 _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7382__S _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4246__S _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5569__C _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4790_ _1617_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__S _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3884__I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5202__I0 _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6460_ _3050_ _2872_ _3052_ _2826_ _3053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_112_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__I0 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5411_ _1905_ memory\[18\]\[2\] _2026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_24_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6391_ _2933_ _2980_ _2984_ _2985_ _2986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5805__S _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8130_ _0430_ clknet_leaf_165_clk_i memory\[26\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5342_ _1957_ memory\[26\]\[1\] _1958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_130_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8061_ _0361_ clknet_leaf_13_clk_i memory\[23\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7012_ memory\[13\]\[15\] _1202_ _3480_ _3486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7091__I _3505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5273_ _1889_ _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4224_ _1299_ _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4155_ _1269_ memory\[15\]\[14\] _1261_ _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6636__S _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5969__A1 _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4086_ _1222_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_104_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7914_ _0214_ clknet_leaf_125_clk_i memory\[1\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4492__I1 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7845_ _0145_ clknet_leaf_142_clk_i memory\[17\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3995__S _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_21_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6371__S _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4988_ memory\[27\]\[10\] _1191_ _1722_ _1723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7776_ _0076_ clknet_leaf_174_clk_i memory\[12\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3939_ net8 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_92_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6727_ _2933_ _3310_ _3312_ _3313_ _3314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__6146__A1 _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7194__I0 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6658_ memory\[20\]\[29\] memory\[21\]\[29\] _1869_ _3246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ _1929_ memory\[11\]\[6\] _2219_ _2174_ _2220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_14_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5942__C _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8328_ _0628_ clknet_leaf_107_clk_i memory\[9\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6589_ memory\[8\]\[27\] memory\[9\]\[27\] _2780_ _3179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6449__A2 _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8259_ _0559_ clknet_leaf_142_clk_i memory\[30\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4180__I0 _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4066__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6281__S _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 data_i[19] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_135_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput27 data_i[29] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_134_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput38 we_i net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5852__C _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6683__C _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5960_ _2515_ memory\[7\]\[13\] _2563_ _2517_ _2564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_88_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5891_ _2163_ _2494_ _2495_ _2496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4911_ _1681_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7287__S _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7630_ memory\[6\]\[17\] net14 _3806_ _3814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4704__S _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_195_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4842_ _1252_ memory\[25\]\[6\] _1638_ _1645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7561_ _3777_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4773_ _1608_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7492_ _3740_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6128__A1 _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6512_ _3101_ _3103_ _2887_ _3104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_132_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6443_ _2000_ memory\[29\]\[24\] _3035_ _2855_ _3036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_15_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6923__I0 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6374_ _2828_ memory\[10\]\[22\] _2969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8113_ _0413_ clknet_leaf_48_clk_i memory\[25\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5325_ _1929_ memory\[2\]\[0\] _1941_ _1942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8044_ _0344_ clknet_leaf_53_clk_i memory\[23\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5639__B1 _2248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5256_ _1872_ _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_110_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4207_ _1302_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5187_ _1114_ memory\[30\]\[8\] _1819_ _1828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_3_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6593__C _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4138_ net37 _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4069_ memory\[12\]\[19\] _1210_ _1192_ _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input19_I data_i[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6603__A2 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7651__I1 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7828_ _0128_ clknet_leaf_33_clk_i memory\[29\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6367__A1 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7759_ _0059_ clknet_leaf_62_clk_i memory\[12\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6119__A1 _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_129_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6276__S _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4524__S _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5581__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4392__I0 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6090_ _2267_ memory\[1\]\[16\] _2690_ _2509_ _2691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5110_ _1787_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7330__I0 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5041_ _1246_ memory\[28\]\[3\] _1747_ _1751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_108_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8731_ _1031_ clknet_leaf_1_clk_i memory\[6\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6992_ _3475_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5943_ memory\[14\]\[13\] _2547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_36_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4434__S _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5874_ _2432_ memory\[26\]\[12\] _2479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_48_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8662_ _0962_ clknet_leaf_206_clk_i memory\[10\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8593_ _0893_ clknet_leaf_69_clk_i memory\[4\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7613_ memory\[6\]\[9\] net37 _3795_ _3805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ _1635_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7544_ _3768_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4756_ net38 _1168_ _1597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7475_ _3731_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4687_ _1559_ _1448_ _1560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_71_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6588__C _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6426_ memory\[2\]\[23\] memory\[3\]\[23\] _2736_ _3020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5492__C _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4383__I0 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6357_ _2754_ _2951_ _2666_ _2952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_8_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5308_ _1879_ _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5999__I _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6288_ memory\[2\]\[20\] memory\[3\]\[20\] _2736_ _2885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_126_Left_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4609__S _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8027_ _0327_ clknet_leaf_39_clk_i memory\[22\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5239_ _1293_ _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7624__I1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6588__A1 _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_212_clk_i clknet_4_0_0_clk_i clknet_leaf_212_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_3_clk_i clknet_4_1_0_clk_i clknet_leaf_3_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_123_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4344__S _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_135_Left_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5239__I _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7655__S _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5683__B _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6760__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5175__S _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6498__C _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3982__I net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7390__S _3686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_143_clk_i_I clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7312__I0 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4519__S _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6019__B _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5251__A1 _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4254__S _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4053__I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_68_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4610_ _1518_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5590_ _1883_ _2199_ _2200_ _2201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4601__I1 _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4541_ _1481_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5085__S _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7260_ _1104_ memory\[3\]\[3\] _3614_ _3618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6503__A1 _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4472_ _1444_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4365__I0 _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6211_ _2754_ _2808_ _2666_ _2809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7191_ _3581_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6142_ _2515_ memory\[7\]\[17\] _2741_ _2517_ _2742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_21_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6909__S _3396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4429__S _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6073_ _1863_ _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4668__I1 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5024_ _1741_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6975_ _1160_ memory\[16\]\[30\] _3432_ _3466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5926_ _2108_ memory\[28\]\[13\] _2530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4164__S _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8714_ _1014_ clknet_leaf_84_clk_i memory\[6\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5487__C _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8645_ _0945_ clknet_leaf_147_clk_i memory\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5857_ _2267_ memory\[1\]\[11\] _2462_ _2043_ _2463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_63_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5788_ memory\[20\]\[10\] memory\[21\]\[10\] _2346_ _2395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4808_ memory\[24\]\[22\] _1217_ _1624_ _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8576_ _0876_ clknet_leaf_170_clk_i memory\[3\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_133_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4739_ _1588_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7527_ memory\[5\]\[0\] net6 _3759_ _3760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7274__I _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7458_ _1093_ memory\[10\]\[0\] _3722_ _3723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4356__I0 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6409_ _2674_ memory\[18\]\[23\] _3003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3859__A2 _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7389_ _3685_ _3686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6819__S _3383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4659__I1 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4138__I net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_151_clk_i clknet_4_10_0_clk_i clknet_leaf_151_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_166_clk_i clknet_4_8_0_clk_i clknet_leaf_166_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_94_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6733__A1 _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5633__S _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_104_clk_i clknet_4_15_0_clk_i clknet_leaf_104_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_119_clk_i clknet_4_14_0_clk_i clknet_leaf_119_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5472__A1 _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6691__C _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3887__I net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6760_ _1905_ memory\[0\]\[31\] _3346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_128_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5711_ _2267_ memory\[1\]\[8\] _2319_ _2043_ _2320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3972_ _1143_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4822__I1 _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6691_ _1903_ memory\[27\]\[30\] _3277_ _1882_ _3278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_58_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8430_ _0730_ clknet_leaf_64_clk_i memory\[13\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5642_ _2208_ memory\[18\]\[7\] _2252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_73_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6724__A1 _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ memory\[4\]\[5\] _1998_ _2185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6212__B _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8361_ _0661_ clknet_leaf_153_clk_i memory\[14\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4524_ memory\[20\]\[20\] _1212_ _1472_ _1473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7312_ _1156_ memory\[3\]\[28\] _3636_ _3645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8292_ _0592_ clknet_leaf_144_clk_i net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7243_ _3608_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4455_ _1068_ memory\[1\]\[20\] _1435_ _1436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5770__C _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4386_ _1068_ memory\[18\]\[20\] _1398_ _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7174_ memory\[11\]\[27\] _1227_ _3564_ _3572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6125_ memory\[12\]\[17\] memory\[13\]\[17\] _2453_ _2725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6056_ _2380_ _2634_ _2656_ _2657_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__3998__S _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5007_ _1732_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_107_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_83_clk_i clknet_4_12_0_clk_i clknet_leaf_83_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_120_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6958_ _3457_ _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ memory\[4\]\[12\] _2468_ _2514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6889_ memory\[14\]\[21\] _1215_ _3419_ _3421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_134_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_98_clk_i clknet_4_13_0_clk_i clknet_leaf_98_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_119_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8628_ _0928_ clknet_leaf_81_clk_i memory\[0\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4622__S _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8559_ _0859_ clknet_leaf_99_clk_i memory\[3\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6122__B _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6191__A2 _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_21_clk_i clknet_4_3_0_clk_i clknet_leaf_21_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_114_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5453__S _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4069__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_16_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5252__I _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_36_clk_i clknet_4_4_0_clk_i clknet_leaf_36_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5454__A1 _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6016__C _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4804__I1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4532__S _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6706__A1 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7506__I0 _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5363__S _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4240_ _1319_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6686__C _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4740__I0 _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6258__I _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4171_ _1239_ _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5445__A1 _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7930_ _0230_ clknet_leaf_208_clk_i memory\[1\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7861_ _0161_ clknet_leaf_26_clk_i memory\[17\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6812_ _1133_ memory\[9\]\[17\] _3372_ _3380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7792_ _0092_ clknet_leaf_62_clk_i memory\[15\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3955_ memory\[19\]\[16\] _1131_ _1119_ _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6743_ memory\[23\]\[31\] _1895_ _3328_ _2006_ _3329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4442__S _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6674_ _1909_ _3261_ _1994_ _3262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_135_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5625_ _1855_ _2214_ _2234_ _2235_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_8413_ _0713_ clknet_leaf_186_clk_i memory\[16\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3886_ _1083_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5337__I _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5556_ _2150_ _2155_ _2159_ _2167_ _1918_ _2168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8344_ _0644_ clknet_leaf_214_clk_i memory\[9\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4507_ memory\[20\]\[12\] _1196_ _1461_ _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8275_ _0575_ clknet_leaf_32_clk_i memory\[30\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5487_ _2084_ _2089_ _2094_ _2100_ _1952_ _2101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4438_ _1265_ memory\[1\]\[12\] _1424_ _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7226_ _3599_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_53_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4369_ _1265_ memory\[18\]\[12\] _1387_ _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7157_ memory\[11\]\[19\] _1210_ _3553_ _3563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6108_ _2529_ memory\[29\]\[17\] _2707_ _2389_ _2708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7088_ _3526_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6039_ _2310_ memory\[11\]\[15\] _2639_ _2640_ _2641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5956__B _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4352__S _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4151__I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6164__A2 _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7663__S _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__I _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5183__S _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5675__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5427__A1 _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6742__S _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4262__S _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7573__S _3781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5902__A2 _2506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6697__B _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5410_ _2022_ _1894_ _2024_ _1901_ _2025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_6390_ _2938_ _2939_ memory\[5\]\[22\] _2985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5341_ _1910_ _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_50_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8060_ _0360_ clknet_leaf_13_clk_i memory\[23\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5093__S _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7011_ _3485_ _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5666__A1 _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5272_ _1165_ _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_10_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4713__I0 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4223_ _1310_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6917__S _3433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_191_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4154_ net11 _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_128_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4085_ memory\[12\]\[24\] _1221_ _1213_ _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5969__A2 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7913_ _0213_ clknet_leaf_111_clk_i memory\[1\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_104_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7844_ _0144_ clknet_leaf_136_clk_i memory\[17\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7775_ _0075_ clknet_leaf_171_clk_i memory\[12\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7547__I _3758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4987_ _1710_ _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_19_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4172__S _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6394__A2 _2964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6726_ _2938_ _2939_ memory\[5\]\[30\] _3313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3938_ _1120_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7483__S _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6146__A2 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6657_ memory\[22\]\[29\] _3245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3869_ net20 _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_33_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5608_ _1930_ memory\[10\]\[6\] _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4900__S _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6588_ _2776_ memory\[11\]\[27\] _3177_ _1907_ _3178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_131_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8327_ _0627_ clknet_leaf_107_clk_i memory\[9\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5539_ _2108_ memory\[28\]\[5\] _2151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4952__I0 _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8258_ _0558_ clknet_leaf_136_clk_i memory\[30\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7209_ _1121_ memory\[8\]\[11\] _3589_ _3591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4704__I0 _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8189_ _0489_ clknet_leaf_4_clk_i memory\[27\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6827__S _3383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5409__B2 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6082__B2 _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7457__I _3721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3985__I net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__A2 _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4082__S _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5906__S _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput17 data_i[1] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput28 data_i[2] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5196__I0 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6688__A3 _3274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4810__S _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5896__B2 _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5705__I _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__B _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6999__I1 _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4056__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5820__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5890_ _1057_ _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_48_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4910_ _1252_ memory\[26\]\[6\] _1674_ _1681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4841_ _1644_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_138_clk_i_I clknet_4_9_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7560_ memory\[5\]\[16\] net13 _3770_ _3777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6204__C _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4772_ memory\[24\]\[5\] _1181_ _1602_ _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7491_ _1131_ memory\[10\]\[16\] _3733_ _3740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_83_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7176__I1 _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6511_ _2884_ _3102_ _1913_ _3103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5187__I0 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6442_ _2001_ memory\[28\]\[24\] _3035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_43_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5887__A1 _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8112_ _0412_ clknet_leaf_48_clk_i memory\[25\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6373_ _2965_ _2872_ _2967_ _2826_ _2968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_100_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5324_ _1882_ _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8043_ _0343_ clknet_leaf_47_clk_i memory\[23\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5639__B2 _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5255_ _1371_ _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6300__A2 _2870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4206_ _1242_ memory\[29\]\[1\] _1300_ _1302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_110_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4167__S _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5186_ _1827_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_3_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4137_ _1257_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7100__I1 _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5111__I0 _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4068_ net16 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_79_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6382__S _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7827_ _0127_ clknet_leaf_33_clk_i memory\[29\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6181__I _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7758_ _0058_ clknet_leaf_63_clk_i memory\[12\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7689_ _3844_ _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6709_ memory\[14\]\[30\] _3296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5953__C _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5327__B1 _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4630__S _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5878__A1 _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4925__I0 _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6055__A1 _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5260__I _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4540__S _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5869__A1 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6905__I1 _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4916__I0 _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5040_ _1750_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6294__A1 _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_64_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5170__I _1818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6991_ memory\[13\]\[5\] _1181_ _3469_ _3475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__S _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5942_ _2528_ _2535_ _2539_ _2545_ _2403_ _2546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_88_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6841__I0 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7298__S _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8730_ _1030_ clknet_leaf_211_clk_i memory\[6\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6597__A2 _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5873_ memory\[24\]\[12\] _2333_ _2478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6349__A2 _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8661_ _0961_ clknet_leaf_203_clk_i memory\[10\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8592_ _0892_ clknet_leaf_67_clk_i memory\[4\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7612_ _3804_ _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4824_ memory\[24\]\[30\] _1233_ _1601_ _1635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7543_ memory\[5\]\[8\] net36 _3759_ _3768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3958__I1 _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4755_ _1596_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7149__I1 _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4450__S _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7474_ _1114_ memory\[10\]\[8\] _3722_ _3731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4686_ net38 _1061_ _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_4_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6425_ _2733_ memory\[1\]\[23\] _3018_ _2975_ _3019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6521__A2 _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6356_ memory\[30\]\[22\] memory\[31\]\[22\] _2532_ _2951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_8_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5307_ memory\[12\]\[0\] memory\[13\]\[0\] _1923_ _1924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8026_ _0326_ clknet_leaf_39_clk_i memory\[22\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5281__S _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6285__A1 _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6287_ _1882_ _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5238_ _1854_ _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input31_I data_i[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6037__A1 _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5169_ _1294_ _1374_ _1818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_98_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5948__C _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3949__I1 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4360__S _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7671__S _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7560__I1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3885__I0 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6823__I0 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4540_ memory\[20\]\[28\] _1229_ _1472_ _1481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_53_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7581__S _3781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4471_ _1084_ memory\[1\]\[28\] _1435_ _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6210_ memory\[30\]\[19\] memory\[31\]\[19\] _2532_ _2808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7190_ _1102_ memory\[8\]\[2\] _3578_ _3581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6141_ _2562_ memory\[6\]\[17\] _2741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6267__A1 _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _2669_ _2294_ _2672_ _2250_ _2673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6925__S _3433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5023_ memory\[27\]\[27\] _1227_ _1733_ _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3876__I0 _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5490__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6814__I0 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6974_ _3465_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8713_ _1013_ clknet_leaf_104_clk_i memory\[6\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5925_ _1861_ _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_75_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5856_ _2318_ memory\[0\]\[11\] _2462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_119_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8644_ _0944_ clknet_leaf_148_clk_i memory\[10\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4807_ _1626_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5787_ memory\[22\]\[10\] _2394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8575_ _0875_ clknet_leaf_168_clk_i memory\[3\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4180__S _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6599__C _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7526_ _3758_ _3759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4738_ _1074_ memory\[23\]\[23\] _1584_ _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4669_ _1550_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7457_ _3721_ _3722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_44_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7491__S _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6408_ _2999_ _2760_ _3001_ _2716_ _3002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_3_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7388_ _1598_ _1411_ _3685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_101_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6339_ memory\[4\]\[21\] _2934_ _2935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8009_ _0309_ clknet_leaf_128_clk_i memory\[22\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6835__S _3383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5481__A2 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3867__I0 _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__C _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6430__A1 _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4154__I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6570__S _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5694__B _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_12_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7230__I0 _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4595__I1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3971_ memory\[19\]\[21\] _1142_ _1140_ _1143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_18_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5710_ _2318_ memory\[0\]\[8\] _2319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_9_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7221__I0 _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6690_ _2898_ memory\[26\]\[30\] _3277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_45_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5641_ _2246_ _1894_ _2249_ _2250_ _2251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_61_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4586__I1 _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5572_ _2181_ _2183_ _1950_ _2184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8360_ _0660_ clknet_leaf_149_clk_i memory\[14\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4523_ _1449_ _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8291_ _0591_ clknet_leaf_140_clk_i net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7311_ _3644_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7242_ _1154_ memory\[8\]\[27\] _3600_ _3608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_2_clk_i clknet_4_0_0_clk_i clknet_leaf_2_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_133_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_211_clk_i clknet_4_0_0_clk_i clknet_leaf_211_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4454_ _1412_ _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4385_ _1375_ _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_55_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7173_ _3571_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6124_ memory\[14\]\[17\] _2724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6055_ _2330_ net45 _2657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5006_ memory\[27\]\[19\] _1210_ _1722_ _1732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_107_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6957_ _1142_ memory\[16\]\[21\] _3455_ _3457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6412__A1 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7460__I0 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4274__I0 _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5908_ _2510_ _2512_ _2421_ _2513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_66_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6888_ _3420_ _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5839_ _2442_ _2294_ _2444_ _2250_ _2445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_118_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8627_ _0927_ clknet_leaf_81_clk_i memory\[0\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6403__B _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_186_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8558_ _0858_ clknet_leaf_98_clk_i memory\[3\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7509_ _3749_ _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8489_ _0789_ clknet_leaf_111_clk_i memory\[11\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5734__S _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7279__I0 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output62_I net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6651__A1 _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3988__I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4085__S _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6403__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7396__S _3686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6032__C _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5644__S _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4170_ _1279_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4059__I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6642__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7690__I0 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7860_ _0160_ clknet_leaf_31_clk_i memory\[17\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6811_ _3379_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7442__I0 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7791_ _0091_ clknet_leaf_62_clk_i memory\[15\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4256__I0 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4723__S _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3954_ net13 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_86_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6742_ memory\[20\]\[31\] memory\[21\]\[31\] _1869_ _3328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6673_ memory\[8\]\[29\] memory\[9\]\[29\] _1992_ _3261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3885_ _1082_ memory\[7\]\[27\] _1066_ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_135_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5624_ _1954_ net67 _2235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8412_ _0712_ clknet_leaf_185_clk_i memory\[16\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4559__I1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8343_ _0643_ clknet_leaf_205_clk_i memory\[9\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5555_ _2162_ _2166_ _1916_ _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_150_clk_i clknet_4_10_0_clk_i clknet_leaf_150_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4506_ _1463_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8274_ _0574_ clknet_leaf_74_clk_i memory\[30\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5486_ _1997_ _2095_ _2098_ _2099_ _2100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_41_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4437_ _1426_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7225_ _1137_ memory\[8\]\[19\] _3589_ _3599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7156_ _3562_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4368_ _1389_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6107_ _2574_ memory\[28\]\[17\] _2707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_165_clk_i clknet_4_8_0_clk_i clknet_leaf_165_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4299_ _1267_ memory\[17\]\[13\] _1347_ _1351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7087_ memory\[31\]\[18\] _1208_ _3517_ _3526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6038_ _1882_ _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_69_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6117__C _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7989_ _0289_ clknet_leaf_37_clk_i memory\[21\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_103_clk_i clknet_4_15_0_clk_i clknet_leaf_103_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6912__I _3432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_118_clk_i clknet_4_11_0_clk_i clknet_leaf_118_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_20_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5263__I _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6321__B1 _2911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5675__A2 _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__S _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6624__B2 _3212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6624__A1 _3198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4789__I1 _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6043__B _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5882__B _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5340_ memory\[24\]\[1\] _1859_ _1956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_130_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_82_clk_i clknet_4_12_0_clk_i clknet_leaf_82_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5271_ _1883_ _1886_ _1887_ _1888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_50_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7010_ memory\[13\]\[14\] _1200_ _3480_ _3485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4222_ _1258_ memory\[29\]\[9\] _1300_ _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_134_clk_i_I clknet_4_9_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4153_ _1268_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_97_clk_i clknet_4_13_0_clk_i clknet_leaf_97_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_128_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7663__I0 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4084_ net22 _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7912_ _0212_ clknet_leaf_112_clk_i memory\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4477__I0 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7415__I0 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4229__I0 _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7843_ _0143_ clknet_leaf_136_clk_i memory\[17\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_20_clk_i clknet_4_3_0_clk_i clknet_leaf_20_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4986_ _1721_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7774_ _0074_ clknet_leaf_169_clk_i memory\[12\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3937_ memory\[19\]\[10\] _1118_ _1119_ _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_63_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6725_ _2981_ memory\[7\]\[30\] _3311_ _2983_ _3312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_clkbuf_leaf_59_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_35_clk_i clknet_4_4_0_clk_i clknet_leaf_35_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6656_ _3241_ _3243_ _1889_ _3244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3868_ _1071_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6587_ _2828_ memory\[10\]\[27\] _3177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5607_ _2215_ _1921_ _2217_ _1927_ _2218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_8326_ _0626_ clknet_leaf_114_clk_i memory\[9\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5538_ _1857_ _2146_ _2148_ _2149_ _2150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_115_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8257_ _0557_ clknet_leaf_134_clk_i memory\[30\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7208_ _3590_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5469_ memory\[15\]\[3\] _1922_ _2082_ _1925_ _2083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_74_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8188_ _0488_ clknet_leaf_6_clk_i memory\[27\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7139_ memory\[11\]\[10\] _1191_ _3553_ _3554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5811__I _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4628__S _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7004__S _3480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5409__A2 _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6606__A1 _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6082__A2 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7406__I0 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 data_i[20] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5194__S _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput29 data_i[30] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5345__A1 _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5896__A2 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5721__I _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4538__S _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4459__I0 _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5596__C _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4840_ _1250_ memory\[25\]\[5\] _1638_ _1644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_60_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6510_ memory\[2\]\[25\] memory\[3\]\[25\] _2736_ _3102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4072__I _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5584__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4771_ _1607_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7490_ _3739_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6441_ _2798_ _3030_ _3032_ _3033_ _3034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_31_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6372_ memory\[15\]\[22\] _2823_ _2966_ _2773_ _2967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8111_ _0411_ clknet_leaf_47_clk_i memory\[25\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5323_ _1933_ _1938_ _1939_ _1940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8042_ _0342_ clknet_leaf_131_clk_i memory\[23\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5639__A2 _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4698__I0 _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5254_ _1870_ _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4448__S _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5185_ _1112_ memory\[30\]\[7\] _1819_ _1827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4205_ _1301_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6300__A3 _2895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4136_ _1256_ memory\[15\]\[8\] _1240_ _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_3_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4067_ _1209_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6663__S _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7826_ _0126_ clknet_leaf_33_clk_i memory\[29\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7757_ _0057_ clknet_leaf_64_clk_i memory\[12\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5575__A1 _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4969_ memory\[27\]\[1\] _1173_ _1711_ _1713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7688_ _1125_ memory\[7\]\[13\] _3837_ _3844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6708_ _3280_ _3285_ _3289_ _3294_ _1094_ _3295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_50_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6639_ memory\[4\]\[28\] _2934_ _3228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4710__I _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8309_ _0609_ clknet_leaf_192_clk_i net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4358__S _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7669__S _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7252__A1 _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4157__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5802__A2 _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4861__I0 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5189__S _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5566__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4268__S _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7579__S _3781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7094__I1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6990_ _3474_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5941_ _2542_ _2544_ _2302_ _2545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5099__S _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5872_ _2380_ _2451_ _2476_ _2477_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_8660_ _0960_ clknet_leaf_80_clk_i memory\[10\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8591_ _0891_ clknet_leaf_67_clk_i memory\[4\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7611_ memory\[6\]\[8\] net36 _3795_ _3804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _1634_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7542_ _3767_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4754_ _1091_ memory\[23\]\[31\] _1561_ _1596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7473_ _3730_ _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5309__B2 _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4685_ _1558_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6424_ _2784_ memory\[0\]\[23\] _3018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_112_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6658__S _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6355_ _2529_ memory\[29\]\[22\] _2949_ _2855_ _2950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_8_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5306_ _1884_ _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6286_ _2733_ memory\[1\]\[20\] _2882_ _2509_ _2883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8025_ _0325_ clknet_leaf_38_clk_i memory\[22\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5237_ net38 _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4178__S _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7489__S _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5168_ _1817_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input24_I data_i[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7085__I1 _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5099_ _1091_ memory\[28\]\[31\] _1746_ _1781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_3_Left_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4906__S _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4119_ _1245_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7809_ _0109_ clknet_leaf_135_clk_i memory\[29\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4641__S _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6899__I1 _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__A1 _2309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4088__S _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_58_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4816__S _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5087__I0 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__I0 _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5539__A1 _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4551__S _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5446__I _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _1443_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5711__A1 _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6140_ memory\[4\]\[17\] _2468_ _2740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6071_ memory\[23\]\[16\] _2247_ _2670_ _2671_ _2672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _1740_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7102__S _3528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5778__A1 _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6973_ _1158_ memory\[16\]\[29\] _3455_ _3465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8712_ _1012_ clknet_leaf_109_clk_i memory\[6\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5924_ _2332_ _2523_ _2525_ _2527_ _2528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_76_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5855_ _2458_ _2460_ _2414_ _2461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_119_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8643_ _0943_ clknet_leaf_149_clk_i memory\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4806_ memory\[24\]\[21\] _1215_ _1624_ _1626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__S _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5786_ _2390_ _2392_ _2291_ _2393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_63_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8574_ _0874_ clknet_leaf_199_clk_i memory\[3\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5950__A1 _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4737_ _1587_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7525_ _3757_ _1485_ _3758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_44_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4668_ memory\[22\]\[23\] _1219_ _1546_ _1550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7456_ _1374_ _3359_ _3721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__5702__A1 _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6407_ memory\[23\]\[23\] _2713_ _3000_ _2671_ _3001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_102_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4599_ memory\[21\]\[23\] _1219_ _1509_ _1513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7387_ _3684_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6338_ _1858_ _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6269_ memory\[16\]\[20\] memory\[17\]\[20\] _2630_ _2866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5466__B1 _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_182_clk_i_I clknet_4_9_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8008_ _0308_ clknet_leaf_121_clk_i memory\[22\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7058__I1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4636__S _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7012__S _3480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6851__S _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5975__B _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4371__S _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6194__A1 _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7682__S _3837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5266__I _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_66_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4546__S _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3970_ net19 _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_75_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5377__S _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5640_ _1058_ _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4035__I1 _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5571_ _1941_ _2182_ _2136_ _2183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ _1471_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8290_ _0590_ clknet_leaf_141_clk_i net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7310_ _1154_ memory\[3\]\[27\] _3636_ _3644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4453_ _1434_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7241_ _3607_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5904__I _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_84_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4384_ _1397_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_55_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7172_ memory\[11\]\[26\] _1225_ _3564_ _3571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6936__S _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6123_ _2706_ _2711_ _2717_ _2722_ _2403_ _2723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_0_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6054_ _2638_ _2645_ _2650_ _2655_ _2428_ _2656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5005_ _1731_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6660__A2 _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_93_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6956_ _3456_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5907_ _2418_ _2511_ _2136_ _2512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_120_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5795__B _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_129_clk_i_I clknet_4_14_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6887_ memory\[14\]\[20\] _1212_ _3419_ _3420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5838_ memory\[23\]\[11\] _2247_ _2443_ _2205_ _2444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8626_ _0926_ clknet_leaf_84_clk_i memory\[0\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4026__I1 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5223__I0 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8557_ _0857_ clknet_4_13_0_clk_i memory\[3\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5923__A1 _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5769_ _1997_ _2373_ _2375_ _2376_ _2377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__6971__I0 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7508_ _1148_ memory\[10\]\[24\] _3744_ _3749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8488_ _0788_ clknet_leaf_114_clk_i memory\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6479__A2 _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5814__I _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7439_ _3712_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6100__A1 _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5750__S _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output55_I net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6380__I _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4017__I1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5914__A1 _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__I _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5599__C _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4276__S _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6642__A2 _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6810_ _1131_ memory\[9\]\[16\] _3372_ _3379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7587__S _3781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4075__I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7790_ _0090_ clknet_leaf_63_clk_i memory\[15\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3953_ _1130_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6741_ memory\[22\]\[31\] _3327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_130_clk_i_I clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__I _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6223__C _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4803__I _1601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6672_ _1987_ memory\[11\]\[29\] _3259_ _1907_ _3260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3884_ net25 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5905__A1 _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5623_ _2218_ _2223_ _2228_ _2233_ _1952_ _2234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_8411_ _0711_ clknet_leaf_185_clk_i memory\[16\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8342_ _0642_ clknet_leaf_204_clk_i memory\[9\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_4_13_0_clk_i clknet_0_clk_i clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5554_ _2163_ _2165_ _2029_ _2166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4505_ memory\[20\]\[11\] _1194_ _1461_ _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8273_ _0573_ clknet_leaf_59_clk_i memory\[30\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5485_ _2005_ _2007_ memory\[5\]\[3\] _2099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4436_ _1263_ memory\[1\]\[11\] _1424_ _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7224_ _3598_ _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6330__A1 _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4367_ _1263_ memory\[18\]\[11\] _1387_ _1389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7155_ memory\[11\]\[18\] _1208_ _3553_ _3562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4192__I0 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5570__S _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6106_ _2332_ _2702_ _2704_ _2705_ _2706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_67_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4298_ _1350_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_55_clk_i_I clknet_4_5_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7086_ _3525_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6037_ _2362_ memory\[10\]\[15\] _2639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4186__S _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5302__C _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7497__S _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4914__S _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7988_ _0288_ clknet_leaf_38_clk_i memory\[21\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6397__A1 _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6939_ _3447_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6149__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8609_ _0909_ clknet_leaf_139_clk_i memory\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6944__I0 _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6308__C _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4486__I1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__S _1601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7200__S _3578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_1_clk_i clknet_4_0_0_clk_i clknet_leaf_1_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_83_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_210_clk_i clknet_4_0_0_clk_i clknet_leaf_210_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7188__I0 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_130_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5270_ _1293_ _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_120_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4221_ _1309_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4174__I0 _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6486__S _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4152_ _1267_ memory\[15\]\[13\] _1261_ _1268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4083_ _1220_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7911_ _0211_ clknet_leaf_113_clk_i memory\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4734__S _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7842_ _0142_ clknet_leaf_137_clk_i memory\[17\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6379__A1 _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7110__S _3528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6234__B _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7773_ _0073_ clknet_leaf_216_clk_i memory\[12\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4985_ memory\[27\]\[9\] _1189_ _1711_ _1721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3936_ _1097_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_63_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6724_ _1864_ memory\[6\]\[30\] _3311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6655_ _1932_ _3242_ _1856_ _3243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3867_ _1070_ memory\[7\]\[21\] _1066_ _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5792__C _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5354__A2 _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6551__A1 _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ _3173_ _2872_ _3175_ _2826_ _3176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5606_ memory\[15\]\[6\] _1922_ _2216_ _1925_ _2217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_103_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8325_ _0625_ clknet_leaf_117_clk_i memory\[9\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5537_ _1871_ _2060_ memory\[25\]\[5\] _2149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_115_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6303__A1 _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8256_ _0556_ clknet_leaf_167_clk_i memory\[2\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7351__I0 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7207_ _1118_ memory\[8\]\[10\] _3589_ _3590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5468_ memory\[12\]\[3\] memory\[13\]\[3\] _1978_ _2082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_74_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4419_ _1246_ memory\[1\]\[3\] _1413_ _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8187_ _0487_ clknet_leaf_6_clk_i memory\[27\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5399_ _1862_ memory\[27\]\[2\] _2013_ _1867_ _2014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_7138_ _3541_ _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7069_ _3516_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_6_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4617__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7020__S _3480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6917__I0 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput19 data_i[21] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_30_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7690__S _3837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6319__B _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7645__I1 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5449__I _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5033__A1 _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_164_clk_i clknet_4_8_0_clk_i clknet_leaf_164_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4770_ memory\[24\]\[4\] _1179_ _1602_ _1607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5584__A2 _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6533__B2 _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6440_ _2803_ _1990_ memory\[25\]\[24\] _3033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_43_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6371_ memory\[12\]\[22\] memory\[13\]\[22\] _2919_ _2966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8110_ _0410_ clknet_leaf_47_clk_i memory\[25\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5322_ _1889_ _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_51_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_179_clk_i clknet_4_8_0_clk_i clknet_leaf_179_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4729__S _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5912__I _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8041_ _0341_ clknet_leaf_130_clk_i memory\[23\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5253_ _1869_ _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_11_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_102_clk_i clknet_4_12_0_clk_i clknet_leaf_102_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5184_ _1826_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4204_ _1237_ memory\[29\]\[0\] _1300_ _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6944__S _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4135_ net36 _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_3_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4066_ memory\[12\]\[18\] _1208_ _1192_ _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_117_clk_i clknet_4_14_0_clk_i clknet_leaf_117_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7825_ _0125_ clknet_leaf_33_clk_i memory\[29\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7756_ _0056_ clknet_leaf_61_clk_i memory\[12\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6772__A1 _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4622__I1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4968_ _1712_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7687_ _3843_ _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3919_ _1107_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6707_ _3291_ _3293_ _1915_ _3294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_50_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5295__S _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4899_ _1675_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5327__A2 _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6638_ _3224_ _3226_ _2887_ _3227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6524__A1 _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4386__I0 _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8308_ _0608_ clknet_leaf_31_clk_i net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6569_ _2000_ memory\[29\]\[27\] _3158_ _2855_ _3159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_14_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7324__I0 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8239_ _0539_ clknet_leaf_97_clk_i memory\[2\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6139__B _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_81_clk_i clknet_4_12_0_clk_i clknet_leaf_81_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4613__I1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6763__A1 _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_177_clk_i_I clknet_4_9_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_96_clk_i clknet_4_13_0_clk_i clknet_leaf_96_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6515__A1 _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4377__I0 _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6321__C _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5933__S _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7618__I1 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_34_clk_i clknet_4_4_0_clk_i clknet_leaf_34_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_18_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4301__I0 _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5940_ _2163_ _2543_ _2495_ _2544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4284__S _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5871_ _2330_ net41 _2477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7610_ _3803_ _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_49_clk_i clknet_4_5_0_clk_i clknet_leaf_49_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7595__S _3795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8590_ _0890_ clknet_leaf_92_clk_i memory\[4\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_60_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4822_ memory\[24\]\[29\] _1231_ _1624_ _1634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7541_ memory\[5\]\[7\] net35 _3759_ _3767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4753_ _1595_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6512__B _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7472_ _1112_ memory\[10\]\[7\] _3722_ _3730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6506__A1 _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5309__A2 _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4684_ memory\[22\]\[31\] _1235_ _1523_ _1558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6423_ _3014_ _3016_ _2880_ _3017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_102_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6354_ _2574_ memory\[28\]\[22\] _2949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7306__I0 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6285_ _2784_ memory\[0\]\[20\] _2882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4459__S _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5305_ _1895_ _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8024_ _0324_ clknet_leaf_38_clk_i memory\[22\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5236_ _1853_ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_71_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5493__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7609__I1 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ _1162_ memory\[2\]\[31\] _1782_ _1817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5098_ _1780_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4118_ _1244_ memory\[15\]\[2\] _1240_ _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4049_ _1197_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input17_I data_i[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4194__S _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6745__A1 _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7808_ _0108_ clknet_leaf_173_clk_i memory\[15\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7739_ _0039_ clknet_leaf_184_clk_i memory\[19\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6422__B _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_104_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6849__S _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5980__C _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4369__S _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5552__I _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5484__A1 _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6584__S _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_113_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6736__A1 _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4832__S _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_122_Left_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_115_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6051__C _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5011__I1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input9_I data_i[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6070_ _1371_ _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_127_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5021_ memory\[27\]\[26\] _1225_ _1733_ _1740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4078__I net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7389__I _3685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6507__B _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8711_ _1011_ clknet_leaf_109_clk_i memory\[6\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6972_ _3464_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5923_ _2337_ _2526_ memory\[25\]\[13\] _2527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5854_ _2313_ _2459_ _2177_ _2460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4742__S _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8642_ _0942_ clknet_leaf_149_clk_i memory\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6727__A1 _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4805_ _1625_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8573_ _0873_ clknet_leaf_199_clk_i memory\[3\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5785_ _2288_ _2391_ _2200_ _2392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7524_ _1057_ _1064_ _3757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5637__I _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4202__A2 _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4736_ _1072_ memory\[23\]\[22\] _1584_ _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5002__I1 _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4667_ _1549_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7455_ _3720_ _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6406_ memory\[20\]\[23\] memory\[21\]\[23\] _2812_ _3000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7386_ _1162_ memory\[4\]\[31\] _3649_ _3684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4598_ _1512_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6337_ _1058_ _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5372__I _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_125_clk_i_I clknet_4_14_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6268_ _2626_ memory\[19\]\[20\] _2864_ _2541_ _2865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5466__A1 _2062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6199_ _2380_ _2770_ _2795_ _2797_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5219_ _1146_ memory\[30\]\[23\] _1841_ _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8007_ _0307_ clknet_leaf_155_clk_i memory\[22\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5321__B _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4816__I1 _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6718__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6194__A2 _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7518__I0 _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6579__S _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4752__I0 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5282__I _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5570_ memory\[2\]\[5\] memory\[3\]\[5\] _1992_ _2182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4521_ memory\[20\]\[19\] _1210_ _1461_ _1471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_123_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4452_ _1056_ memory\[1\]\[19\] _1424_ _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3906__S _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7240_ _1152_ memory\[8\]\[26\] _3600_ _3607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5406__B _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4383_ _1056_ memory\[18\]\[19\] _1387_ _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_55_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7171_ _3570_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6122_ _2719_ _2721_ _2302_ _2722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5448__A1 _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6053_ _2467_ _2651_ _2653_ _2654_ _2655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5004_ memory\[27\]\[18\] _1208_ _1722_ _1731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_37_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6952__S _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6955_ _1139_ memory\[16\]\[20\] _3455_ _3456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5906_ memory\[2\]\[12\] memory\[3\]\[12\] _2270_ _2511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_120_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5620__A1 _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8625_ _0925_ clknet_leaf_100_clk_i memory\[0\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_66_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6886_ _3396_ _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_134_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5837_ memory\[20\]\[11\] memory\[21\]\[11\] _2346_ _2443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_51_clk_i_I clknet_4_5_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6176__A2 _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4271__I _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8556_ _0856_ clknet_leaf_105_clk_i memory\[3\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5923__A2 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5768_ _2005_ _2007_ memory\[5\]\[9\] _2376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4719_ _1269_ memory\[23\]\[14\] _1573_ _1578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8487_ _0787_ clknet_leaf_116_clk_i memory\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7507_ _3748_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5699_ memory\[15\]\[8\] _1922_ _2306_ _2307_ _2308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7438_ _1146_ memory\[0\]\[23\] _3708_ _3712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5687__B2 _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4734__I0 _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7369_ _3675_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4647__S _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5439__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7023__S _3491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output48_I net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5611__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5478__S _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5277__I _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5914__A2 _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7116__A1 _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__A1 _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4725__I0 _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4557__S _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6627__B1 _3215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6740_ _3323_ _3325_ _1889_ _3326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_133_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3952_ memory\[19\]\[15\] _1129_ _1119_ _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6504__C _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6671_ _1988_ memory\[10\]\[29\] _3259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3883_ _1081_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_135_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5622_ _1997_ _2229_ _2231_ _2232_ _2233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_8410_ _0710_ clknet_leaf_188_clk_i memory\[16\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5553_ memory\[16\]\[5\] memory\[17\]\[5\] _2164_ _2165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8341_ _0641_ clknet_leaf_200_clk_i memory\[9\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _1462_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7108__S _3528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8272_ _0572_ clknet_leaf_61_clk_i memory\[30\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5669__A1 _2261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5484_ _2049_ memory\[7\]\[3\] _2097_ _2051_ _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4435_ _1425_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7223_ _1135_ memory\[8\]\[18\] _3589_ _3598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7154_ _3561_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4366_ _1388_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6105_ _2337_ _2526_ memory\[25\]\[17\] _2705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_10_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4467__S _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4297_ _1265_ memory\[17\]\[12\] _1347_ _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7130__I1 _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7085_ memory\[31\]\[17\] _1206_ _3517_ _3525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6036_ _2635_ _2406_ _2637_ _2360_ _2638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__5841__A1 _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7987_ _0287_ clknet_leaf_42_clk_i memory\[21\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6938_ _1123_ memory\[16\]\[12\] _3444_ _3447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6414__C _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6869_ _3410_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8608_ _0908_ clknet_leaf_175_clk_i memory\[4\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8539_ _0839_ clknet_leaf_213_clk_i memory\[8\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7018__S _3480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__S _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4377__S _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6085__A1 _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3930__I1 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5132__I0 _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__A1 _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7688__S _3837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4840__S _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5899__A1 _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4946__I0 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4220_ _1256_ memory\[29\]\[8\] _1300_ _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4151_ net10 _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3921__I1 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7112__I1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5403__C _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4082_ memory\[12\]\[23\] _1219_ _1213_ _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5823__A1 _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7910_ _0210_ clknet_leaf_113_clk_i memory\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7841_ _0141_ clknet_leaf_137_clk_i memory\[17\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7772_ _0072_ clknet_leaf_218_clk_i memory\[12\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4984_ _1720_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3935_ net7 _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_74_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6723_ memory\[4\]\[30\] _2934_ _3310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4750__S _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6654_ memory\[30\]\[29\] memory\[31\]\[29\] _1923_ _3242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6000__A1 _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3866_ net19 _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5605_ memory\[12\]\[6\] memory\[13\]\[6\] _1978_ _2216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4937__I0 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6585_ memory\[15\]\[27\] _2823_ _3174_ _2773_ _3175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_27_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8324_ _0624_ clknet_leaf_118_clk_i memory\[9\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5536_ _1862_ memory\[27\]\[5\] _2147_ _1867_ _2148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_115_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8255_ _0555_ clknet_leaf_168_clk_i memory\[2\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5467_ memory\[14\]\[3\] _2081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_112_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7206_ _3577_ _3589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4418_ _1416_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8186_ _0486_ clknet_leaf_4_clk_i memory\[27\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5398_ _1957_ memory\[26\]\[2\] _2013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7137_ _3552_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_74_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3912__I1 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4349_ _1379_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7068_ memory\[31\]\[9\] _1189_ _3506_ _3516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6019_ _2618_ _2620_ _2291_ _2621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4925__S _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6058__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6386__I _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_173_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5290__I _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5105__I0 _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7211__S _3589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6335__B _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6054__C _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5893__C _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_98_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4919__I0 _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6533__A2 _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7581__I1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6370_ memory\[14\]\[22\] _2965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5321_ _1934_ _1936_ _1937_ _1938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8040_ _0340_ clknet_leaf_121_clk_i memory\[23\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5252_ _1059_ _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5183_ _1110_ memory\[30\]\[6\] _1819_ _1826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4203_ _1299_ _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_110_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6229__C _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4134_ _1255_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_3_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4065_ net15 _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_79_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7824_ _0124_ clknet_leaf_56_clk_i memory\[29\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6221__A1 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7755_ _0055_ clknet_leaf_77_clk_i memory\[12\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4967_ memory\[27\]\[0\] _1164_ _1711_ _1712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7686_ _1123_ memory\[7\]\[12\] _3837_ _3843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_62_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3918_ memory\[19\]\[4\] _1106_ _1098_ _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6706_ _1873_ _3292_ _2961_ _3293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_50_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4898_ _1237_ memory\[26\]\[0\] _1674_ _1675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_105_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6524__A2 _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6637_ _2884_ _3225_ _1913_ _3226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_105_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6568_ _2001_ memory\[28\]\[27\] _3158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_132_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8307_ _0607_ clknet_leaf_32_clk_i net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5519_ _2129_ _2131_ _1939_ _2132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_76_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6499_ memory\[14\]\[25\] _3091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_0_clk_i clknet_4_0_0_clk_i clknet_leaf_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8238_ _0538_ clknet_leaf_105_clk_i memory\[2\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8169_ _0469_ clknet_leaf_176_clk_i memory\[27\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4655__S _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6835__I0 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7031__S _3491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6870__S _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4454__I _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5994__B _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7260__I0 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4390__S _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6763__A2 _3348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6602__C _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6279__A1 _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3888__I0 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5888__C _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4565__S _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6844__I _3396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6451__A1 _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5870_ _2456_ _2461_ _2466_ _2475_ _2428_ _2476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__4364__I _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6203__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4821_ _1633_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7675__I _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6754__A2 _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3909__S _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7540_ _3766_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4752_ _1089_ memory\[23\]\[30\] _1561_ _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_60_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7471_ _3729_ _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4683_ _1557_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7554__I1 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6422_ _2779_ _3015_ _2643_ _3016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6353_ _2798_ _2944_ _2946_ _2947_ _2948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_11_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6284_ _2877_ _2879_ _2880_ _2881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5304_ _1893_ _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_110_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8023_ _0323_ clknet_leaf_38_clk_i memory\[22\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6955__S _3455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5235_ _1162_ memory\[30\]\[31\] _1818_ _1853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_71_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6690__A1 _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3879__I0 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5493__A2 _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4540__I1 _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5166_ _1816_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4117_ net28 _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5097_ _1089_ memory\[28\]\[30\] _1746_ _1780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4475__S _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4048_ memory\[12\]\[12\] _1196_ _1192_ _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6442__A1 _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7242__I0 _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5999_ _1238_ _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_leaf_121_clk_i_I clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7807_ _0107_ clknet_leaf_172_clk_i memory\[15\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4756__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7738_ _0038_ clknet_leaf_189_clk_i memory\[19\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7545__I1 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7669_ _1106_ memory\[7\]\[4\] _1087_ _3834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_62_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6808__I0 _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_46_clk_i_I clknet_4_5_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_163_clk_i clknet_4_10_0_clk_i clknet_leaf_163_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7481__I0 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6433__A1 _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4295__I0 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7696__S _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_178_clk_i clknet_4_9_0_clk_i clknet_leaf_178_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_85_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6613__B _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_101_clk_i clknet_4_13_0_clk_i clknet_leaf_101_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5944__S _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_116_clk_i clknet_4_14_0_clk_i clknet_leaf_116_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4770__I1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5020_ _1739_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6672__A1 _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4295__S _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7472__I0 _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6424__A1 _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4286__I0 _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8710_ _1010_ clknet_leaf_108_clk_i memory\[6\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6971_ _1156_ memory\[16\]\[28\] _3455_ _3464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5922_ _1872_ _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5853_ memory\[8\]\[11\] memory\[9\]\[11\] _2314_ _2459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8641_ _0941_ clknet_leaf_149_clk_i memory\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5784_ memory\[30\]\[10\] memory\[31\]\[10\] _2066_ _2391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4804_ memory\[24\]\[20\] _1212_ _1624_ _1625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8572_ _0872_ clknet_leaf_201_clk_i memory\[3\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4735_ _1586_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7523_ _3756_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ memory\[22\]\[22\] _1217_ _1546_ _1549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7454_ _1162_ memory\[0\]\[31\] _3685_ _3720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4597_ memory\[21\]\[22\] _1217_ _1509_ _1512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6405_ memory\[22\]\[23\] _2999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4210__I0 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7385_ _3683_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6336_ _2929_ _2931_ _2887_ _2932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xclkbuf_leaf_80_clk_i clknet_4_6_0_clk_i clknet_leaf_80_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_110_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6267_ _2674_ memory\[18\]\[20\] _2864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4513__I1 _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6198_ _2796_ net48 _2797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5218_ _1844_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8006_ _0306_ clknet_leaf_161_clk_i memory\[22\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5602__B _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3901__I _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5149_ _1144_ memory\[2\]\[22\] _1805_ _1808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_95_clk_i clknet_4_13_0_clk_i clknet_leaf_95_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7215__I0 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4933__S _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_33_clk_i clknet_4_4_0_clk_i clknet_leaf_33_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_90_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_48_clk_i clknet_4_5_0_clk_i clknet_leaf_48_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5004__S _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7454__I0 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5939__S _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4268__I0 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8557__CLK clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5738__I _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4440__I0 _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5393__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4520_ _1470_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4451_ _1433_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7170_ memory\[11\]\[25\] _1223_ _3564_ _3570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6121_ _2629_ _2720_ _2495_ _2721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4382_ _1396_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_55_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6052_ _2472_ _2473_ memory\[5\]\[15\] _2654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6645__A1 _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5003_ _1730_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6237__C _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6954_ _3432_ _3455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5905_ _2267_ memory\[1\]\[12\] _2508_ _2509_ _2510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_120_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8624_ _0924_ clknet_leaf_96_clk_i memory\[0\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6885_ _3418_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_66_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5836_ memory\[22\]\[11\] _2442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8555_ _0855_ clknet_leaf_110_clk_i memory\[3\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4431__I0 _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5767_ _2049_ memory\[7\]\[9\] _2374_ _2051_ _2375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_8_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4718_ _1577_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8486_ _0786_ clknet_leaf_116_clk_i memory\[11\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7506_ _1146_ memory\[10\]\[23\] _3744_ _3748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5698_ _1879_ _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4649_ memory\[22\]\[14\] _1200_ _1535_ _1540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7437_ _3711_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5687__A2 _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7368_ _1144_ memory\[4\]\[22\] _3672_ _3675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5316__C _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6319_ _2629_ _2914_ _2495_ _2915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7304__S _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7299_ _3638_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_219_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7684__I0 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5332__B _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6428__B _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7436__I0 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5986__C _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5375__A1 _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4973__I1 _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5293__I _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4838__S _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6627__B2 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7427__I0 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5850__A2 _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3951_ net12 _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_129_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3882_ _1080_ memory\[7\]\[26\] _1066_ _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6670_ _3255_ _2872_ _3257_ _1901_ _3258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_5621_ _2005_ _2007_ memory\[5\]\[6\] _2232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4413__I0 _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_168_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5366__A1 _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8340_ _0640_ clknet_leaf_80_clk_i memory\[9\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5552_ _1884_ _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_5_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8271_ _0571_ clknet_leaf_59_clk_i memory\[30\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4503_ memory\[20\]\[10\] _1191_ _1461_ _1462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5483_ _2096_ memory\[6\]\[3\] _2097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_41_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7222_ _3597_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_117_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4434_ _1260_ memory\[1\]\[10\] _1424_ _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7153_ memory\[11\]\[17\] _1206_ _3553_ _3561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4365_ _1260_ memory\[18\]\[10\] _1387_ _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4748__S _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_220_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7084_ _3524_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6104_ _2382_ memory\[27\]\[17\] _2703_ _2384_ _2704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7124__S _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6035_ memory\[15\]\[15\] _2357_ _2636_ _2307_ _2637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_4296_ _1349_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6094__A2 _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6963__S _3455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7986_ _0286_ clknet_leaf_44_clk_i memory\[21\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6937_ _3446_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5378__I _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6868_ memory\[14\]\[11\] _1194_ _3408_ _3410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_7_0_clk_i clknet_0_clk_i clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_107_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5819_ _2005_ _2007_ memory\[5\]\[10\] _2426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_106_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4404__I0 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8607_ _0907_ clknet_leaf_187_clk_i memory\[4\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6799_ _3373_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8538_ _0838_ clknet_leaf_205_clk_i memory\[8\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8469_ _0769_ clknet_leaf_19_clk_i memory\[31\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6609__A1 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output60_I net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6880__I1 _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5288__I _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7209__S _3589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5520__A1 _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4150_ _1266_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_52_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_94_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6783__S _3361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4081_ net21 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_37_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5823__A2 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7840_ _0140_ clknet_leaf_181_clk_i memory\[29\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4882__I0 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6515__C _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5587__A1 _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7771_ _0071_ clknet_leaf_217_clk_i memory\[12\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4983_ memory\[27\]\[8\] _1187_ _1711_ _1720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3934_ _1117_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_63_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6722_ _3306_ _3308_ _1916_ _3309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6653_ _2000_ memory\[29\]\[29\] _3240_ _2855_ _3241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5339__A1 _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3865_ _1069_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5604_ memory\[14\]\[6\] _2215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6584_ memory\[12\]\[27\] memory\[13\]\[27\] _2919_ _3174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8323_ _0623_ clknet_leaf_118_clk_i memory\[9\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5535_ _1957_ memory\[26\]\[5\] _2147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5466_ _2062_ _2069_ _2073_ _2079_ _1918_ _2080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_8254_ _0554_ clknet_leaf_169_clk_i memory\[2\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7205_ _3588_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4417_ _1244_ memory\[1\]\[2\] _1413_ _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8185_ _0485_ clknet_leaf_9_clk_i memory\[27\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5397_ memory\[24\]\[2\] _1859_ _2012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7136_ memory\[11\]\[9\] _1189_ _3542_ _3552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_74_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4348_ _1244_ memory\[18\]\[2\] _1376_ _1379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7067_ _3515_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4279_ _1340_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6018_ _2288_ _2619_ _2200_ _2620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6706__B _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6425__C _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5578__A1 _2172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7969_ _0269_ clknet_leaf_167_clk_i memory\[21\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7029__S _3491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6868__S _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4388__S _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_116_clk_i_I clknet_4_14_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5504__C _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6853__I1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5569__A1 _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4851__S _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5041__I0 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5320_ _1238_ _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5251_ _1862_ memory\[27\]\[0\] _1865_ _1867_ _1868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4202_ _1294_ _1298_ _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_48_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ _1825_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6049__A2 _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4133_ _1254_ memory\[15\]\[7\] _1240_ _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7402__S _3686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3930__S _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4064_ _1207_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4855__I0 _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7823_ _0123_ clknet_leaf_46_clk_i memory\[29\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_125_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7754_ _0054_ clknet_leaf_178_clk_i memory\[12\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6705_ memory\[16\]\[30\] memory\[17\]\[30\] _1885_ _3292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4966_ _1710_ _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_19_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7685_ _3842_ _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3917_ net32 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6261__B _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4897_ _1673_ _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_105_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6636_ memory\[2\]\[28\] memory\[3\]\[28\] _1911_ _3225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5732__A1 _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6567_ _2798_ _3153_ _3155_ _3156_ _3157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_113_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8306_ _0606_ clknet_leaf_73_clk_i net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5518_ _1934_ _2130_ _1937_ _2131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_76_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6498_ _3075_ _3080_ _3084_ _3089_ _2869_ _3090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_8237_ _0537_ clknet_leaf_98_clk_i memory\[2\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5449_ _1861_ _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5391__I _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4001__S _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8168_ _0468_ clknet_leaf_139_clk_i memory\[27\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7119_ _3543_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5099__I0 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7312__S _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8099_ _0399_ clknet_leaf_175_clk_i memory\[25\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4846__I0 _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6460__A2 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_42_clk_i_I clknet_4_4_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7012__I1 _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5723__A1 _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7079__I1 _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4846__S _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4820_ memory\[24\]\[28\] _1229_ _1624_ _1633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5962__A1 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4751_ _1594_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_60_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7470_ _1110_ memory\[10\]\[6\] _3722_ _3729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4682_ memory\[22\]\[30\] _1233_ _1523_ _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6421_ memory\[8\]\[23\] memory\[9\]\[23\] _2780_ _3015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6352_ _2803_ _2526_ memory\[25\]\[22\] _2947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_59_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5425__B _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6283_ _1889_ _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5303_ memory\[14\]\[0\] _1920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8022_ _0322_ clknet_leaf_37_clk_i memory\[22\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5234_ _1852_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5165_ _1160_ memory\[2\]\[30\] _1782_ _1816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7132__S _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4116_ _1243_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5096_ _1779_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4047_ net9 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6971__S _3455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7806_ _0106_ clknet_leaf_171_clk_i memory\[15\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5998_ memory\[2\]\[14\] memory\[3\]\[14\] _2270_ _2601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5953__A1 _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7737_ _0037_ clknet_leaf_20_clk_i memory\[19\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4949_ _1701_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7668_ _3833_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6619_ _1877_ memory\[18\]\[28\] _3208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7599_ memory\[6\]\[2\] net28 _3795_ _3798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_18_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4666__S _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6681__A2 _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_27_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5296__I _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7217__S _3589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_123_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6121__A1 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4576__S _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5899__C _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6791__S _3361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6970_ _3463_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5921_ _2382_ memory\[27\]\[13\] _2524_ _2384_ _2525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_109_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5200__S _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5852_ _2310_ memory\[11\]\[11\] _2457_ _2174_ _2458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_119_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5235__I0 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6523__C _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8640_ _0940_ clknet_leaf_174_clk_i memory\[0\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4038__I1 _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5783_ _2063_ memory\[29\]\[10\] _2388_ _2389_ _2390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_75_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4803_ _1601_ _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8571_ _0871_ clknet_leaf_204_clk_i memory\[3\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_32_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4734_ _1070_ memory\[23\]\[21\] _1584_ _1586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7522_ _1162_ memory\[10\]\[31\] _3721_ _3756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4665_ _1548_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_54_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7453_ _3719_ _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4596_ _1511_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6404_ _2995_ _2997_ _2757_ _2998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7384_ _1160_ memory\[4\]\[30\] _3649_ _3683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6335_ _2884_ _2930_ _2602_ _2931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6266_ _2860_ _2760_ _2862_ _2716_ _2863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8005_ _0305_ clknet_leaf_162_clk_i memory\[22\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6197_ _1854_ _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5217_ _1144_ memory\[30\]\[22\] _1841_ _1844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4486__S _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5148_ _1807_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input22_I data_i[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5079_ _1070_ memory\[28\]\[21\] _1769_ _1771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_84_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6179__A1 _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_215_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4029__I1 _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5926__A1 _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_2_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_10_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7037__S _3491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6351__A1 _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6876__S _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6103__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4396__S _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7500__S _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_18_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5217__I0 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5917__A1 _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6965__I0 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6590__A1 _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5754__I _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4450_ _1277_ memory\[1\]\[18\] _1424_ _1433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7390__I0 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4381_ _1277_ memory\[18\]\[18\] _1387_ _1396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_133_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6120_ memory\[16\]\[17\] memory\[17\]\[17\] _2630_ _2720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_55_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _2515_ memory\[7\]\[15\] _2652_ _2517_ _2653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_56_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6645__A2 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5002_ memory\[27\]\[17\] _1206_ _1722_ _1730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_164_clk_i_I clknet_4_8_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6518__C _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6953_ _3454_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_120_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5208__I0 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6884_ memory\[14\]\[19\] _1210_ _3408_ _3418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5904_ _1879_ _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8623_ _0923_ clknet_leaf_99_clk_i memory\[0\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5835_ _2438_ _2440_ _2291_ _2441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_66_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8554_ _0854_ clknet_leaf_88_clk_i memory\[3\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5766_ _2096_ memory\[6\]\[9\] _2374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_62_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_162_clk_i clknet_4_10_0_clk_i clknet_leaf_162_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_127_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4717_ _1267_ memory\[23\]\[13\] _1573_ _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_89_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8485_ _0785_ clknet_leaf_147_clk_i memory\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7505_ _3747_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5697_ memory\[12\]\[8\] memory\[13\]\[8\] _1978_ _2306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4648_ _1539_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7436_ _1144_ memory\[0\]\[22\] _3708_ _3711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6333__A1 _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6696__S _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4579_ _1502_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7367_ _3674_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_177_clk_i clknet_4_9_0_clk_i clknet_leaf_177_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6318_ memory\[16\]\[21\] memory\[17\]\[21\] _2630_ _2914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7298_ _1142_ memory\[3\]\[21\] _3636_ _3638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_3_0_clk_i clknet_0_clk_i clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6249_ _1854_ _2846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_100_clk_i clknet_4_13_0_clk_i clknet_leaf_100_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4498__I1 _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5105__S _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4944__S _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_115_clk_i clknet_4_15_0_clk_i clknet_leaf_115_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4670__I1 _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7372__I0 _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4186__I0 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4918__I _1673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6627__A2 _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5015__S _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7230__S _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5749__I _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3950_ _1128_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6938__I0 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3881_ net24 _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5620_ _2049_ memory\[7\]\[6\] _2230_ _2051_ _2231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_42_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_90_clk_i_I clknet_4_13_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5551_ _1872_ _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8270_ _0570_ clknet_leaf_60_clk_i memory\[30\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4502_ _1449_ _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5417__C _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7221_ _1133_ memory\[8\]\[17\] _3589_ _3597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_94_clk_i clknet_4_13_0_clk_i clknet_leaf_94_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_111_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5482_ _1863_ _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_117_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3933__S _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4433_ _1412_ _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_1_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7152_ _3560_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4364_ _1375_ _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6529__B _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7083_ memory\[31\]\[16\] _1204_ _3517_ _3524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4295_ _1263_ memory\[17\]\[11\] _1347_ _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6079__B1 _2673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6103_ _2432_ memory\[26\]\[17\] _2703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6618__A2 _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6034_ memory\[12\]\[15\] memory\[13\]\[15\] _2453_ _2636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_32_clk_i clknet_4_6_0_clk_i clknet_leaf_32_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_68_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4764__S _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7985_ _0285_ clknet_leaf_50_clk_i memory\[21\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6936_ _1121_ memory\[16\]\[11\] _3444_ _3446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_47_clk_i clknet_4_5_0_clk_i clknet_leaf_47_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6867_ _3409_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6929__I0 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6798_ _1118_ memory\[9\]\[10\] _3372_ _3373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5818_ _2049_ memory\[7\]\[10\] _2424_ _2051_ _2425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8606_ _0906_ clknet_leaf_172_clk_i memory\[4\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5749_ _1895_ _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_8_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8537_ _0837_ clknet_leaf_205_clk_i memory\[8\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6306__A1 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8468_ _0768_ clknet_leaf_30_clk_i memory\[31\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7419_ _1127_ memory\[0\]\[14\] _3697_ _3702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8399_ _0699_ clknet_leaf_100_clk_i memory\[16\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7657__I1 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output53_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5997__C _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4674__S _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7050__S _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4643__I1 _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5596__A2 _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_112_clk_i_I clknet_4_15_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A1 _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5518__B _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7345__I0 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7225__S _3589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_52_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_37_clk_i_I clknet_4_4_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4080_ _1218_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4584__S _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5700__C _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4634__I1 _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4982_ _1719_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7770_ _0070_ clknet_leaf_216_clk_i memory\[12\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3933_ memory\[19\]\[9\] _1116_ _1098_ _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6721_ _1883_ _3307_ _1913_ _3308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6652_ _2001_ memory\[28\]\[29\] _3240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6536__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3864_ _1068_ memory\[7\]\[20\] _1066_ _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5603_ _2196_ _2202_ _2207_ _2213_ _1918_ _2214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4398__I0 _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8322_ _0622_ clknet_leaf_146_clk_i memory\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6583_ memory\[14\]\[27\] _3173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7336__I0 _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5534_ memory\[24\]\[5\] _1859_ _2146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5465_ _2076_ _2078_ _1916_ _2079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8253_ _0553_ clknet_leaf_200_clk_i memory\[2\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7204_ _1116_ memory\[8\]\[9\] _3578_ _3588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8184_ _0484_ clknet_leaf_10_clk_i memory\[27\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4416_ _1415_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7135_ _3551_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5396_ _1855_ _1976_ _2010_ _2011_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__7639__I1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4347_ _1378_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7066_ memory\[31\]\[8\] _1187_ _3506_ _3515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4278_ _1246_ memory\[17\]\[3\] _1336_ _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6017_ memory\[30\]\[15\] memory\[31\]\[15\] _2532_ _2619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4322__I0 _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4494__S _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5389__I _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7968_ _0268_ clknet_leaf_131_clk_i memory\[20\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6775__A1 _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7899_ _0199_ clknet_leaf_25_clk_i memory\[18\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6919_ _1104_ memory\[16\]\[3\] _3433_ _3437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6722__B _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6527__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__S _3468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6884__S _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5299__I _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6766__A1 _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6632__B _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6351__C _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5741__A2 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7318__I0 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5250_ _1866_ _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_121_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ _1297_ _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5181_ _1108_ memory\[30\]\[5\] _1819_ _1825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4132_ net35 _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4063_ memory\[12\]\[17\] _1206_ _1192_ _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5257__A1 _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7822_ _0122_ clknet_leaf_57_clk_i memory\[29\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4607__I1 _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4965_ _1709_ _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_47_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7753_ _0053_ clknet_leaf_154_clk_i memory\[12\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6034__S _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5937__I _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3916_ _1105_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6704_ _1876_ memory\[19\]\[30\] _3290_ _2003_ _3291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6509__A1 _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5980__A2 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7684_ _1121_ memory\[7\]\[11\] _3837_ _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4896_ _1374_ _1599_ _1673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_50_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6635_ _1904_ memory\[1\]\[28\] _3223_ _2975_ _3224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6969__S _3455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6566_ _2803_ _1990_ memory\[25\]\[27\] _3156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_6_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8305_ _0605_ clknet_leaf_58_clk_i net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5517_ memory\[8\]\[4\] memory\[9\]\[4\] _1935_ _2130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_76_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8236_ _0536_ clknet_leaf_105_clk_i memory\[2\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6497_ _3086_ _3088_ _2768_ _3089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_100_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5496__A1 _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5448_ _1857_ _2057_ _2059_ _2061_ _2062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_100_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5379_ _1941_ _1993_ _1994_ _1995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8167_ _0467_ clknet_leaf_155_clk_i memory\[27\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7118_ memory\[11\]\[0\] _1164_ _3542_ _3543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8098_ _0398_ clknet_leaf_175_clk_i memory\[25\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7049_ _3505_ _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5248__A1 _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6717__B _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3920__I net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5113__S _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__A1 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4952__S _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__I _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5420__B2 _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6171__C _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5023__I1 _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5487__A1 _2084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4198__I _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6346__C _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5023__S _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_clk_i_I clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6739__A1 _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__I _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5411__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4750_ _1086_ memory\[23\]\[29\] _1584_ _1594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_60_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6789__S _3361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4681_ _1556_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6420_ _2776_ memory\[11\]\[23\] _3013_ _2640_ _3014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6351_ _2848_ memory\[27\]\[22\] _2945_ _2850_ _2946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_52_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5302_ _1875_ _1891_ _1902_ _1917_ _1918_ _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6282_ _2779_ _2878_ _2643_ _2879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8021_ _0321_ clknet_leaf_36_clk_i memory\[22\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5233_ _1160_ memory\[30\]\[30\] _1818_ _1852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7413__S _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5164_ _1815_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4115_ _1242_ memory\[15\]\[1\] _1240_ _1243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6029__S _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5095_ _1086_ memory\[28\]\[29\] _1769_ _1779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4046_ _1195_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__S _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5650__B2 _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7805_ _0105_ clknet_leaf_194_clk_i memory\[15\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5997_ _2267_ memory\[1\]\[14\] _2599_ _2509_ _2600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4571__I _1486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5402__A1 _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7736_ _0036_ clknet_leaf_25_clk_i memory\[19\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4948_ _1076_ memory\[26\]\[24\] _1696_ _1701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_6_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7667_ _1104_ memory\[7\]\[3\] _1087_ _3833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4879_ _1664_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_159_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6618_ _3204_ _1893_ _3206_ _1937_ _3207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_46_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5616__B _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7598_ _3797_ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6549_ _3137_ _3139_ _2880_ _3140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_30_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8219_ _0519_ clknet_leaf_8_clk_i memory\[28\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5469__B2 _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_211_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6166__C _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4682__S _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_133_Right_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4481__I _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6402__S _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6201__I _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4857__S _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__B _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5920_ _2432_ memory\[26\]\[13\] _2524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_109_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__A1 _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ _2362_ memory\[10\]\[11\] _2457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6092__B _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5935__A2 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5782_ _1879_ _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4802_ _1623_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8570_ _0870_ clknet_leaf_204_clk_i memory\[3\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_32_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4733_ _1585_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_160_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6983__I1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7521_ _3755_ _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7408__S _3686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7452_ _1160_ memory\[0\]\[30\] _3685_ _3719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4664_ memory\[22\]\[21\] _1215_ _1546_ _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6403_ _2754_ _2996_ _2666_ _2997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5699__B2 _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4595_ memory\[21\]\[21\] _1215_ _1509_ _1511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4746__I0 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7383_ _3682_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6334_ memory\[2\]\[21\] memory\[3\]\[21\] _2736_ _2930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6265_ memory\[23\]\[20\] _2713_ _2861_ _2671_ _2862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__7143__S _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5171__I0 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5216_ _1843_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7160__I1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8004_ _0304_ clknet_leaf_161_clk_i memory\[22\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5871__A1 _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6196_ _2775_ _2783_ _2789_ _2794_ _2428_ _2795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5147_ _1142_ memory\[2\]\[21\] _1805_ _1807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_85_clk_i_I clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5078_ _1770_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input15_I data_i[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5623__A1 _2218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4029_ memory\[12\]\[6\] _1183_ _1171_ _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_84_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6714__C _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7719_ _0019_ clknet_leaf_123_clk_i memory\[19\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7318__S _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8699_ _0999_ clknet_leaf_0_clk_i memory\[5\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_4_6_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7117__I _3541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7151__I1 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5614__A1 _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6624__C _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5917__A2 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7228__S _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4380_ _1395_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6087__B _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_107_clk_i_I clknet_4_15_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6050_ _2562_ memory\[6\]\[15\] _2652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5703__C _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5302__B1 _1902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__I0 _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input7_I data_i[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ _1729_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_0_Left_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4900__I0 _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6952_ _1137_ memory\[16\]\[19\] _3444_ _3454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6534__C _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5903_ _2318_ memory\[0\]\[12\] _2508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6883_ _3417_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8622_ _0922_ clknet_leaf_99_clk_i memory\[0\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5834_ _2288_ _2439_ _2200_ _2440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_66_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6030__A1 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8553_ _0853_ clknet_leaf_111_clk_i memory\[3\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5765_ memory\[4\]\[9\] _1998_ _2373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4716_ _1576_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8484_ _0784_ clknet_leaf_148_clk_i memory\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5696_ memory\[14\]\[8\] _2305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7504_ _1144_ memory\[10\]\[22\] _3744_ _3747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4719__I0 _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4647_ memory\[22\]\[13\] _1198_ _1535_ _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6977__S _3432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7435_ _3710_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7366_ _1142_ memory\[4\]\[21\] _3672_ _3674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4578_ memory\[21\]\[13\] _1198_ _1498_ _1502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_102_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6776__I _3360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6317_ _2626_ memory\[19\]\[21\] _2912_ _2541_ _2913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_12_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6097__A1 _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7297_ _3637_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6248_ _2380_ _2821_ _2844_ _2845_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6179_ _2776_ memory\[11\]\[18\] _2777_ _2640_ _2778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_99_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7601__S _3795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5121__S _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4960__S _1673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4958__I0 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6887__S _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3933__I1 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7124__I1 _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5031__S _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6012__A1 _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3880_ _1079_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6563__A2 _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_33_clk_i_I clknet_4_4_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5550_ _2160_ memory\[19\]\[5\] _2161_ _2075_ _2162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_5_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4501_ _1460_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5481_ memory\[4\]\[3\] _1998_ _2095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7220_ _3596_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4432_ _1423_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6315__A2 _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7151_ memory\[11\]\[16\] _1204_ _3553_ _3560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5714__B _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5206__S _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4363_ _1386_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3924__I1 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7082_ _3523_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5126__I0 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4294_ _1348_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6102_ memory\[24\]\[17\] _2333_ _2702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6033_ memory\[14\]\[15\] _2635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7421__S _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7984_ _0284_ clknet_leaf_50_clk_i memory\[21\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6935_ _3445_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4780__S _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6003__A1 _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6866_ memory\[14\]\[10\] _1191_ _3408_ _3409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5817_ _2096_ memory\[6\]\[10\] _2424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6797_ _3360_ _3372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8605_ _0905_ clknet_leaf_194_clk_i memory\[4\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5748_ memory\[14\]\[9\] _2356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8536_ _0836_ clknet_leaf_214_clk_i memory\[8\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8467_ _0767_ clknet_leaf_32_clk_i memory\[31\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5679_ _1882_ _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_79_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6500__S _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7418_ _3701_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8398_ _0698_ clknet_leaf_103_clk_i memory\[16\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7349_ _1125_ memory\[4\]\[13\] _3661_ _3665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3923__I net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3915__I1 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7106__I1 _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5117__I0 _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6439__C _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4020__S _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5343__C _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5817__A1 _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6455__B _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6242__A1 _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4690__S _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6190__B _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7506__S _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_81_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_130_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3906__I1 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput70 net70 data_o[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_52_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4865__S _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6481__A1 _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_161_clk_i clknet_4_10_0_clk_i clknet_leaf_161_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_90_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_47_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7281__I0 _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ memory\[27\]\[7\] _1185_ _1711_ _1719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3932_ net37 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_86_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6720_ memory\[2\]\[30\] memory\[3\]\[30\] _1911_ _3307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_176_clk_i clknet_4_8_0_clk_i clknet_leaf_176_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_129_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5495__I _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6651_ _1887_ _3235_ _3237_ _3238_ _3239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_46_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3863_ net18 _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_119_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5602_ _2210_ _2212_ _1916_ _2213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6582_ _3157_ _3162_ _3166_ _3171_ _2869_ _3172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_15_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5533_ _1855_ _2123_ _2144_ _2145_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_8321_ _0621_ clknet_leaf_147_clk_i memory\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5464_ _1909_ _2077_ _2029_ _2078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8252_ _0552_ clknet_leaf_199_clk_i memory\[2\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7203_ _3587_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_114_clk_i clknet_4_15_0_clk_i clknet_leaf_114_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8183_ _0483_ clknet_leaf_10_clk_i memory\[27\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4415_ _1242_ memory\[1\]\[1\] _1413_ _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5395_ _1954_ net50 _2011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7134_ memory\[11\]\[8\] _1187_ _3542_ _3551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6259__C _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4346_ _1242_ memory\[18\]\[1\] _1376_ _1378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7151__S _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7065_ _3514_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4277_ _1339_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_129_Left_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6016_ _2529_ memory\[29\]\[15\] _2617_ _2389_ _2618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_leaf_129_clk_i clknet_4_14_0_clk_i clknet_leaf_129_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6472__A1 _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7272__I0 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7967_ _0267_ clknet_leaf_132_clk_i memory\[20\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7898_ _0198_ clknet_leaf_25_clk_i memory\[18\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6918_ _3436_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_25_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6849_ memory\[14\]\[2\] _1175_ _3397_ _3400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7575__I1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8519_ _0819_ clknet_leaf_107_clk_i memory\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7326__S _3650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4561__I1 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_93_clk_i clknet_4_13_0_clk_i clknet_leaf_93_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_206_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7566__I1 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7236__S _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_31_clk_i clknet_4_6_0_clk_i clknet_leaf_31_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6079__C _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4200_ net38 _1296_ _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_46_clk_i clknet_4_5_0_clk_i clknet_leaf_46_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5180_ _1824_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6829__I0 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4595__S _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4131_ _1253_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5711__C _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4062_ net14 _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6454__A1 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5257__A2 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6206__A1 _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7254__I0 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7821_ _0121_ clknet_leaf_57_clk_i memory\[29\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4964_ _1062_ _1599_ _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_59_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7752_ _0052_ clknet_leaf_150_clk_i memory\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3915_ memory\[19\]\[3\] _1104_ _1098_ _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6703_ _1877_ memory\[18\]\[30\] _3290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_129_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7683_ _3841_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4895_ _1672_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6634_ _1905_ memory\[0\]\[28\] _3223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_73_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6565_ _2848_ memory\[27\]\[27\] _3154_ _2850_ _3155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_6_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8304_ _0604_ clknet_leaf_59_clk_i net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4791__I1 _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5516_ _1929_ memory\[11\]\[4\] _2128_ _1932_ _2129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_6496_ _1873_ _3087_ _2961_ _3088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8235_ _0535_ clknet_leaf_103_clk_i memory\[2\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6985__S _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5447_ _1871_ _2060_ memory\[25\]\[3\] _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_112_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6693__A1 _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5378_ _1238_ _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8166_ _0466_ clknet_leaf_156_clk_i memory\[27\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5902__B _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7117_ _3541_ _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4329_ _1366_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8097_ _0397_ clknet_leaf_175_clk_i memory\[25\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_2_clk_i_I clknet_4_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7493__I0 _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7048_ _3504_ _3505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6445__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_155_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4759__A1 _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5349__B _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6452__C _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5420__A2 _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7548__I1 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6024__I _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4231__I0 _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5723__A3 _2329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7056__S _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6895__S _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6684__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4534__I1 _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5531__C _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7236__I0 _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6362__C _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5974__S _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7539__I1 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4680_ memory\[22\]\[29\] _1231_ _1546_ _1556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5773__I _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4222__I0 _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6350_ _2898_ memory\[26\]\[22\] _2945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6911__A2 _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5301_ _1094_ _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_110_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6281_ memory\[8\]\[20\] memory\[9\]\[20\] _2780_ _2878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_110_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8020_ _0320_ clknet_leaf_34_clk_i memory\[22\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5232_ _1851_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5163_ _1158_ memory\[2\]\[29\] _1805_ _1815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4114_ net17 _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6427__A1 _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5094_ _1778_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4045_ memory\[12\]\[11\] _1194_ _1192_ _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6553__B _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5650__A2 _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7804_ _0104_ clknet_leaf_0_clk_i memory\[15\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5996_ _2318_ memory\[0\]\[14\] _2599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_35_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5884__S _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7735_ _0035_ clknet_leaf_24_clk_i memory\[19\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4947_ _1700_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4461__I0 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7666_ _3832_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4878_ _1074_ memory\[25\]\[23\] _1660_ _1664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_81_clk_i_I clknet_4_12_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6617_ memory\[23\]\[28\] _1895_ _3205_ _2006_ _3206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_132_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7597_ memory\[6\]\[1\] net17 _3795_ _3797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6548_ _2779_ _3138_ _1994_ _3139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4764__I1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6479_ memory\[24\]\[25\] _2799_ _3071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8218_ _0518_ clknet_leaf_12_clk_i memory\[28\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6666__B2 _3253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5469__A2 _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8149_ _0449_ clknet_leaf_36_clk_i memory\[26\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5124__S _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7466__I0 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5641__A2 _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4452__I0 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4204__I0 _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7514__S _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4507__I1 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5542__B _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6638__B _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6409__A1 _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7209__I0 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5850_ _2452_ _2406_ _2455_ _2360_ _2456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_122_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5781_ _2108_ memory\[28\]\[10\] _2388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4801_ memory\[24\]\[19\] _1210_ _1613_ _1623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4199__A2 _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5396__A1 _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_103_clk_i_I clknet_4_15_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4994__I1 _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4732_ _1068_ memory\[23\]\[20\] _1584_ _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7520_ _1160_ memory\[10\]\[30\] _3721_ _3755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4663_ _1547_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7451_ _3718_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6402_ memory\[30\]\[23\] memory\[31\]\[23\] _1923_ _2996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5699__A2 _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4594_ _1510_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7382_ _1158_ memory\[4\]\[29\] _3672_ _3682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3952__S _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5008__I _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6333_ _2733_ memory\[1\]\[21\] _2928_ _2509_ _2929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_110_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7696__I0 _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6264_ memory\[20\]\[20\] memory\[21\]\[20\] _2812_ _2861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6648__A1 _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5215_ _1142_ memory\[30\]\[21\] _1841_ _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6548__B _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8003_ _0303_ clknet_leaf_166_clk_i memory\[22\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6195_ _2467_ _2790_ _2792_ _2793_ _2794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__7448__I0 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_13_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_28_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5146_ _1806_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4783__S _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5077_ _1068_ memory\[28\]\[20\] _1769_ _1770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4028_ net34 _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_84_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5979_ memory\[23\]\[14\] _2247_ _2581_ _2205_ _2582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4434__I0 _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7718_ _0018_ clknet_leaf_122_clk_i memory\[19\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4985__I1 _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8698_ _0998_ clknet_leaf_211_clk_i memory\[5\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3926__I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5119__S _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6302__I _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4023__S _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7649_ memory\[6\]\[26\] net24 _3817_ _3824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4958__S _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7334__S _3650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4425__I0 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5029__S _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5550__A1 _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7678__I0 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7244__S _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6368__B _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5000_ memory\[27\]\[16\] _1204_ _1722_ _1729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6951_ _3453_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5902_ _2504_ _2506_ _2414_ _2507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6882_ memory\[14\]\[18\] _1208_ _3408_ _3417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8621_ _0921_ clknet_leaf_99_clk_i memory\[0\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5833_ memory\[30\]\[11\] memory\[31\]\[11\] _2066_ _2439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5369__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7419__S _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8552_ _0852_ clknet_leaf_110_clk_i memory\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_101_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5764_ _2369_ _2371_ _1950_ _2372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_84_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7503_ _3746_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4967__I1 _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4715_ _1265_ memory\[23\]\[12\] _1573_ _1576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5695_ _2285_ _2292_ _2297_ _2303_ _1918_ _2304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_8483_ _0783_ clknet_leaf_148_clk_i memory\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4646_ _1538_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7434_ _1142_ memory\[0\]\[21\] _3708_ _3710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4577_ _1501_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4778__S _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7365_ _3673_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7669__I0 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6316_ _2674_ memory\[18\]\[21\] _2912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6097__A2 _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7296_ _1139_ memory\[3\]\[20\] _3636_ _3637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6247_ _2796_ net49 _2845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6993__S _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_110_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6178_ _2362_ memory\[10\]\[18\] _2777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3855__A1 _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5129_ _1797_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6725__C _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6233__S _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__C _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5780__A1 _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5532__A1 _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7064__S _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5804__C _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4894__I0 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6635__C _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5599__A1 _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7060__I1 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5771__A1 _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4500_ memory\[20\]\[9\] _1189_ _1450_ _1460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5480_ _2091_ _2093_ _1950_ _2094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4431_ _1258_ memory\[1\]\[9\] _1413_ _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_117_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7150_ _3559_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4362_ _1258_ memory\[18\]\[9\] _1376_ _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7081_ memory\[31\]\[15\] _1202_ _3517_ _3523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6101_ _2380_ _2680_ _2700_ _2701_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4293_ _1260_ memory\[17\]\[10\] _1347_ _1348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6874__I1 _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6032_ _2616_ _2621_ _2625_ _2633_ _2403_ _2634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6318__S _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7983_ _0283_ clknet_leaf_51_clk_i memory\[21\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_68_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6934_ _1118_ memory\[16\]\[10\] _3444_ _3445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7149__S _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _3396_ _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8604_ _0904_ clknet_leaf_18_clk_i memory\[4\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5062__I0 _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6796_ _3371_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5816_ memory\[4\]\[10\] _1998_ _2423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6280__C _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5747_ _2339_ _2344_ _2349_ _2354_ _1918_ _2355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_45_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8535_ _0835_ clknet_leaf_206_clk_i memory\[8\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8466_ _0766_ clknet_leaf_33_clk_i memory\[31\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7417_ _1125_ memory\[0\]\[13\] _3697_ _3701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5678_ _2063_ memory\[29\]\[8\] _2286_ _1880_ _2287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_79_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8397_ _0697_ clknet_leaf_101_clk_i memory\[16\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4629_ _1529_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4301__S _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7348_ _3664_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_92_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7279_ _1123_ memory\[3\]\[12\] _3625_ _3628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4876__I0 _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5132__S _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6027__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4971__S _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5866__I _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5053__I0 _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5815__B _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5505__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5307__S _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_128_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_52_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput60 net60 data_o[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_clkbuf_leaf_202_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7522__S _3721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4010__I _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4867__I0 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7321__I _3649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4980_ _1718_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5992__A1 _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3931_ _1115_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3862_ _1067_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_63_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6650_ _1870_ _1990_ memory\[25\]\[29\] _3238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7033__I1 _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5601_ _2163_ _2211_ _2029_ _2212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6581_ _3168_ _3170_ _2768_ _3171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_39_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5532_ _1954_ net65 _2145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8320_ _0620_ clknet_leaf_178_clk_i net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5463_ memory\[16\]\[3\] memory\[17\]\[3\] _1911_ _2077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5217__S _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8251_ _0551_ clknet_leaf_201_clk_i memory\[2\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7202_ _1114_ memory\[8\]\[8\] _3578_ _3587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8182_ _0482_ clknet_leaf_11_clk_i memory\[27\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4414_ _1414_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5394_ _1981_ _1986_ _1996_ _2009_ _1952_ _2010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_41_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4121__S _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7133_ _3550_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4345_ _1377_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7432__S _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6847__I1 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7064_ memory\[31\]\[7\] _1185_ _3506_ _3514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4276_ _1244_ memory\[17\]\[2\] _1336_ _1339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6015_ _2574_ memory\[28\]\[15\] _2617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4791__S _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7966_ _0266_ clknet_leaf_30_clk_i memory\[20\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7897_ _0197_ clknet_leaf_21_clk_i memory\[18\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6917_ _1102_ memory\[16\]\[2\] _3433_ _3436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_25_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6291__B _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5035__I0 _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6848_ _3399_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5735__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_151_clk_i_I clknet_4_10_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7607__S _3795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8518_ _0818_ clknet_leaf_115_clk_i memory\[8\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6783__I0 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ _1100_ memory\[9\]\[1\] _3361_ _3363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5635__B _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8449_ _0749_ clknet_leaf_134_clk_i memory\[31\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5354__C _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3870__S _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5370__B _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_76_clk_i_I clknet_4_6_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6980__I _3468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4206__S _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6421__S _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5037__S _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6151__A1 _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5264__C _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4876__S _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4001__I1 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4130_ _1252_ memory\[15\]\[6\] _1240_ _1253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4061_ _1205_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7820_ _0120_ clknet_leaf_57_clk_i memory\[29\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6206__A2 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5965__A1 _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4963_ _1708_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7751_ _0051_ clknet_leaf_158_clk_i memory\[12\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7006__I1 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7682_ _1118_ memory\[7\]\[10\] _3837_ _3841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3914_ net31 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6702_ _3286_ _1893_ _3288_ _1937_ _3289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_59_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5717__A1 _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4894_ _1091_ memory\[25\]\[31\] _1637_ _1672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_62_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6633_ _3219_ _3221_ _2880_ _3222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_7_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3955__S _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7427__S _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6564_ _2898_ memory\[26\]\[27\] _3154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6390__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8303_ _0603_ clknet_leaf_57_clk_i net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5455__B _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5515_ _1930_ memory\[10\]\[4\] _2128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6495_ memory\[16\]\[25\] memory\[17\]\[25\] _1885_ _3087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6142__A1 _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8234_ _0534_ clknet_leaf_88_clk_i memory\[2\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5446_ _2006_ _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7190__I0 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5377_ memory\[2\]\[1\] memory\[3\]\[1\] _1992_ _1993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7162__S _3564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8165_ _0465_ clknet_leaf_163_clk_i memory\[27\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7116_ _1238_ _1559_ _3358_ _3541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_8096_ _0396_ clknet_leaf_133_clk_i memory\[24\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4328_ _1082_ memory\[17\]\[27\] _1358_ _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input38_I we_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7047_ _1062_ _1294_ _3504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4259_ _1329_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6733__C _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7949_ _0249_ clknet_leaf_53_clk_i memory\[20\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3929__I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4026__S _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6381__A1 _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_160_clk_i clknet_4_10_0_clk_i clknet_leaf_160_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_131_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4696__S _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6684__A2 _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_175_clk_i clknet_4_8_0_clk_i clknet_leaf_175_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6436__A2 _3008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6416__S _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5947__A1 _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_113_clk_i clknet_4_14_0_clk_i clknet_leaf_113_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_128_clk_i clknet_4_14_0_clk_i clknet_leaf_128_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_52_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6372__B2 _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ _1908_ _1914_ _1916_ _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6280_ _2776_ memory\[11\]\[20\] _2876_ _2640_ _2877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_121_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4686__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5231_ _1158_ memory\[30\]\[29\] _1841_ _1851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_71_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5162_ _1814_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5093_ _1084_ memory\[28\]\[28\] _1769_ _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6427__A2 _3020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4113_ _1241_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4044_ net8 _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5938__A1 _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7803_ _0103_ clknet_leaf_217_clk_i memory\[15\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5995_ _2595_ _2597_ _2414_ _2598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_91_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7734_ _0034_ clknet_leaf_24_clk_i memory\[19\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4946_ _1074_ memory\[26\]\[23\] _1696_ _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7157__S _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7665_ _1102_ memory\[7\]\[2\] _1087_ _3832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4877_ _1663_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6616_ memory\[20\]\[28\] memory\[21\]\[28\] _2812_ _3205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7596_ _3796_ _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_24_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6363__A1 _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6547_ memory\[8\]\[26\] memory\[9\]\[26\] _2780_ _3138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_92_clk_i clknet_4_13_0_clk_i clknet_leaf_92_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6115__B2 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6478_ _2846_ _3049_ _3069_ _3070_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_8217_ _0517_ clknet_leaf_13_clk_i memory\[28\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5429_ _1987_ memory\[1\]\[2\] _2042_ _2043_ _2044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8148_ _0448_ clknet_leaf_34_clk_i memory\[26\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5632__C _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6728__C _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6418__A2 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8079_ _0379_ clknet_leaf_50_clk_i memory\[24\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7620__S _3806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5140__S _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_30_clk_i clknet_4_6_0_clk_i clknet_leaf_30_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5229__I0 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6977__I0 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_45_clk_i clknet_4_5_0_clk_i clknet_leaf_45_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6354__A1 _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6106__A1 _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_109_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6373__C _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4800_ _1622_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5780_ _2332_ _2381_ _2385_ _2386_ _2387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_56_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6593__A1 _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4731_ _1561_ _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_29_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5717__C _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4662_ memory\[22\]\[20\] _1212_ _1546_ _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7450_ _1158_ memory\[0\]\[29\] _3708_ _3718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6345__A1 _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6401_ _2000_ memory\[29\]\[23\] _2994_ _2855_ _2995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_198_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4593_ memory\[21\]\[20\] _1212_ _1509_ _1510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7381_ _3681_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6332_ _2784_ memory\[0\]\[21\] _2928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_122_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6263_ memory\[22\]\[20\] _2860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_23_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5214_ _1842_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8002_ _0302_ clknet_leaf_165_clk_i memory\[22\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5225__S _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6194_ _2472_ _2473_ memory\[5\]\[18\] _2793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_86_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5145_ _1139_ memory\[2\]\[20\] _1805_ _1806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7440__S _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5076_ _1746_ _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4027_ _1182_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_84_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4682__I1 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5895__S _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6959__I0 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5978_ memory\[20\]\[14\] memory\[21\]\[14\] _2346_ _2581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7620__I1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5908__B _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4929_ _1271_ memory\[26\]\[15\] _1685_ _1691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7717_ _0017_ clknet_leaf_143_clk_i memory\[19\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8697_ _0997_ clknet_leaf_1_clk_i memory\[5\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7648_ _3823_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7384__I0 _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7579_ memory\[5\]\[25\] net23 _3781_ _3787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6739__B _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3942__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6639__A2 _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output69_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5311__A2 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6193__C _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7611__I1 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6575__B2 _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4214__S _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6327__A1 _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5045__S _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3852__I _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4884__S _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7260__S _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6384__B _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6950_ _1135_ memory\[16\]\[18\] _3444_ _3453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5901_ _2313_ _2505_ _2177_ _2506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_88_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4664__I1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6881_ _3416_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8620_ _0920_ clknet_leaf_104_clk_i memory\[0\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5832_ _2063_ memory\[29\]\[11\] _2437_ _2389_ _2438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_66_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6566__A1 _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8551_ _0851_ clknet_leaf_114_clk_i memory\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5763_ _1941_ _2370_ _2136_ _2371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4714_ _1575_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7502_ _1142_ memory\[10\]\[21\] _3744_ _3746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4124__S _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5694_ _2299_ _2301_ _2302_ _2303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8482_ _0782_ clknet_leaf_148_clk_i memory\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7366__I0 _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4645_ memory\[22\]\[12\] _1196_ _1535_ _1538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7433_ _3709_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4576_ memory\[21\]\[12\] _1196_ _1498_ _1501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_130_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7364_ _1139_ memory\[4\]\[20\] _3672_ _3673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6315_ _2908_ _2760_ _2910_ _2716_ _2911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_12_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7295_ _3613_ _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6278__C _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6246_ _2827_ _2833_ _2838_ _2843_ _2428_ _2844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6177_ _1903_ _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4352__I0 _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7170__S _3564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5128_ _1265_ memory\[2\]\[12\] _1794_ _1797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3855__A2 _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input20_I data_i[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5059_ _1760_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4655__I1 _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6557__A1 _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8749_ _1049_ clknet_leaf_92_clk_i memory\[7\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7357__I0 _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7345__S _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4969__S _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3873__S _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6469__B _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_146_clk_i_I clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6548__A1 _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_135_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5771__A2 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4430_ _1422_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6100_ _2330_ net46 _2701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4361_ _1385_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7080_ _3522_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4292_ _1335_ _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_10_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7520__I0 _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6031_ _2628_ _2632_ _2302_ _2633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4334__I0 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7982_ _0282_ clknet_leaf_52_clk_i memory\[21\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6933_ _3432_ _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_119_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3958__S _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6864_ _3407_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6334__S _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5815_ _2417_ _2420_ _2421_ _2422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_92_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8603_ _0903_ clknet_leaf_209_clk_i memory\[4\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6795_ _1116_ memory\[9\]\[9\] _3361_ _3371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6133__I _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5746_ _2351_ _2353_ _2302_ _2354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8534_ _0834_ clknet_leaf_205_clk_i memory\[8\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8465_ _0765_ clknet_leaf_59_clk_i memory\[31\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4789__S _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5677_ _2108_ memory\[28\]\[8\] _2286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5905__C _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7416_ _3700_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_79_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4628_ memory\[22\]\[4\] _1179_ _1524_ _1529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8396_ _0696_ clknet_leaf_104_clk_i memory\[16\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5514__A2 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6289__B _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6711__B2 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7347_ _1123_ memory\[4\]\[12\] _3661_ _3664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_92_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4559_ memory\[21\]\[4\] _1179_ _1487_ _1492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7278_ _3627_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6229_ _2822_ _2406_ _2825_ _2826_ _2827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__5413__S _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5212__I _1818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4628__I1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4029__S _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5450__A1 _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4005__A2 _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5753__A2 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_72_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7075__S _3517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput50 net50 data_o[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput61 net61 data_o[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7502__I0 _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4316__I0 _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5550__C _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6769__A1 _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3930_ memory\[19\]\[8\] _1114_ _1098_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5441__A1 _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6381__C _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5993__S _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7049__I _3505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3861_ _1056_ memory\[7\]\[19\] _1066_ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5600_ memory\[16\]\[6\] memory\[17\]\[6\] _2164_ _2211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6580_ _1873_ _3169_ _2961_ _3170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5531_ _2127_ _2132_ _2138_ _2143_ _1952_ _2144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_42_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4402__S _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8250_ _0550_ clknet_leaf_203_clk_i memory\[2\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7201_ _3586_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5462_ _1904_ memory\[19\]\[3\] _2074_ _2075_ _2076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_78_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5393_ _1997_ _1999_ _2004_ _2008_ _2009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_8181_ _0481_ clknet_leaf_13_clk_i memory\[27\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4413_ _1237_ memory\[1\]\[0\] _1413_ _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7132_ memory\[11\]\[7\] _1185_ _3542_ _3550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4344_ _1237_ memory\[18\]\[0\] _1376_ _1377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4307__I0 _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7063_ _3513_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_74_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__S _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6014_ _2332_ _2612_ _2614_ _2615_ _2616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4275_ _1338_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5233__S _1818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_6_Left_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6064__S _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7965_ _0265_ clknet_leaf_37_clk_i memory\[20\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4871__I _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6572__B _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7896_ _0196_ clknet_leaf_29_clk_i memory\[18\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6916_ _3435_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6847_ memory\[14\]\[1\] _1173_ _3397_ _3399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6999__S _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6778_ _3362_ _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8517_ _0817_ clknet_leaf_117_clk_i memory\[8\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5729_ _1870_ _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_18_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5408__S _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5499__A1 _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8448_ _0748_ clknet_leaf_173_clk_i memory\[13\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8379_ _0679_ clknet_leaf_0_clk_i memory\[14\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4111__I _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_19_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output51_I net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5671__A1 _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6038__I _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5423__A1 _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5726__A2 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4222__S _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6151__A2 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7533__S _3759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5053__S _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3860__I _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4060_ memory\[12\]\[16\] _1204_ _1192_ _1205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5988__S _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5662__A1 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4892__S _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4962_ _1091_ memory\[26\]\[31\] _1673_ _1708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7750_ _0050_ clknet_leaf_159_clk_i memory\[12\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7681_ _3840_ _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6701_ memory\[23\]\[30\] _1895_ _3287_ _2006_ _3288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4893_ _1671_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3913_ _1103_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_104_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6632_ _1909_ _3220_ _1994_ _3221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6612__S _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5017__I1 _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5736__B _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6563_ memory\[24\]\[27\] _2799_ _3153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6390__A2 _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8302_ _0602_ clknet_leaf_59_clk_i net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6494_ _1876_ memory\[19\]\[25\] _3085_ _2003_ _3086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_30_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5514_ _2124_ _1921_ _2126_ _1927_ _2127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_124_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8233_ _0533_ clknet_leaf_110_clk_i memory\[2\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5445_ _1862_ memory\[27\]\[3\] _2058_ _1867_ _2059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__3971__S _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8164_ _0464_ clknet_leaf_163_clk_i memory\[27\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5376_ _1910_ _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7115_ _3540_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8095_ _0395_ clknet_leaf_183_clk_i memory\[24\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4327_ _1365_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6286__C _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_20_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4258_ _1080_ memory\[29\]\[26\] _1322_ _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7046_ _3503_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5653__A1 _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4700__I0 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4189_ _1289_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_87_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5405__A1 _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6602__B1 _3186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7948_ _0248_ clknet_leaf_52_clk_i memory\[20\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4307__S _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7618__S _3806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7879_ _0179_ clknet_leaf_125_clk_i memory\[18\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5646__B _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3945__I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5138__S _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4042__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5365__C _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4977__S _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7353__S _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5192__I0 _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6196__C _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_69_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6995__I1 _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_78_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6372__A2 _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5230_ _1850_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7172__I1 _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5183__I0 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4686__A2 _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_87_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5161_ _1156_ memory\[2\]\[28\] _1805_ _1814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_71_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5092_ _1777_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4112_ _1237_ memory\[15\]\[0\] _1240_ _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4043_ _1193_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_194_clk_i_I clknet_4_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7388__A1 _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5994_ _2313_ _2596_ _2177_ _2597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4127__S _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7802_ _0102_ clknet_leaf_217_clk_i memory\[15\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_220_clk_i clknet_4_0_0_clk_i clknet_leaf_220_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5310__I _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6060__A1 _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7733_ _0033_ clknet_leaf_25_clk_i memory\[19\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4945_ _1699_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_96_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7438__S _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4876_ _1072_ memory\[25\]\[22\] _1660_ _1663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7664_ _3831_ _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6615_ memory\[22\]\[28\] _3204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7595_ memory\[6\]\[0\] net6 _3795_ _3796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6546_ _2776_ memory\[11\]\[26\] _3136_ _1907_ _3137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4797__S _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6115__A2 _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6477_ _2796_ net55 _3070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5913__C _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8216_ _0516_ clknet_leaf_13_clk_i memory\[28\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5428_ _1872_ _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5874__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4921__I0 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8147_ _0447_ clknet_leaf_44_clk_i memory\[26\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5359_ _1972_ _1974_ _1916_ _1975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8078_ _0378_ clknet_leaf_54_clk_i memory\[24\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7029_ memory\[13\]\[23\] _1219_ _3491_ _3495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6744__C _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6051__A1 _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3876__S _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7083__S _3517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5890__I _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4500__S _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5165__I0 _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6901__I1 _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6000__B _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5865__A1 _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4912__I0 _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5331__S _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6042__A1 _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7258__S _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4730_ _1583_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6162__S _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4661_ _1523_ _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_43_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6400_ _2574_ memory\[28\]\[23\] _2994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_43_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7380_ _1156_ memory\[4\]\[28\] _3672_ _3681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4592_ _1486_ _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6331_ _2924_ _2926_ _2880_ _2927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_24_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7145__I1 _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5733__C _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6262_ _2856_ _2858_ _2757_ _2859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_12_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5856__A1 _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6193_ _2515_ memory\[7\]\[18\] _2791_ _2517_ _2792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_86_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5213_ _1139_ memory\[30\]\[20\] _1841_ _1842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8001_ _0301_ clknet_leaf_165_clk_i memory\[22\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5144_ _1782_ _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_20_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5305__I _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5608__A1 _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5075_ _1768_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4026_ memory\[12\]\[5\] _1181_ _1171_ _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6136__I _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ memory\[22\]\[14\] _2580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7168__S _3564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6580__B _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4928_ _1690_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7716_ _0016_ clknet_leaf_142_clk_i memory\[19\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_174_clk_i clknet_4_8_0_clk_i clknet_leaf_174_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8696_ _0996_ clknet_leaf_1_clk_i memory\[5\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7647_ memory\[6\]\[25\] net23 _3817_ _3823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6800__S _3372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4859_ _1269_ memory\[25\]\[14\] _1649_ _1654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_189_clk_i clknet_4_3_0_clk_i clknet_leaf_189_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7578_ _3786_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7136__I1 _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6529_ _2754_ _3119_ _1856_ _3120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5643__C _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4320__S _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5147__I0 _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_112_clk_i clknet_4_15_0_clk_i clknet_leaf_112_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_31_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5151__S _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_127_clk_i clknet_4_12_0_clk_i clknet_leaf_127_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4990__S _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6575__A2 _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5818__C _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_142_clk_i_I clknet_4_11_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7524__A1 _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6710__S _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__B _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5138__I0 _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6649__C _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5838__B2 _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7541__S _3759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6665__B _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_67_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5900_ memory\[8\]\[12\] memory\[9\]\[12\] _2314_ _2505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6015__A1 _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_91_clk_i clknet_4_13_0_clk_i clknet_leaf_91_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6880_ memory\[14\]\[17\] _1206_ _3408_ _3416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_17_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5831_ _2108_ memory\[28\]\[11\] _2437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6566__A2 _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6810__I0 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5762_ memory\[2\]\[9\] memory\[3\]\[9\] _2270_ _2370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8550_ _0850_ clknet_leaf_116_clk_i memory\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_66_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5728__C _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4713_ _1263_ memory\[23\]\[11\] _1573_ _1575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7501_ _3745_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5693_ _1915_ _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_60_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8481_ _0781_ clknet_leaf_149_clk_i memory\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4644_ _1537_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7432_ _1139_ memory\[0\]\[20\] _3708_ _3709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4575_ _1500_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3927__I1 _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7118__I1 _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7363_ _3649_ _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7294_ _3635_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6314_ memory\[23\]\[21\] _2713_ _2909_ _2671_ _2910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5829__A1 _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6245_ _2467_ _2839_ _2841_ _2842_ _2843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_110_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_44_clk_i clknet_4_4_0_clk_i clknet_leaf_44_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6176_ _2771_ _2406_ _2774_ _2360_ _2775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5127_ _1796_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_137_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5058_ _1263_ memory\[28\]\[11\] _1758_ _1760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6254__A1 _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6294__C _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input13_I data_i[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4009_ _1167_ _1169_ _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xclkbuf_leaf_59_clk_i clknet_4_7_0_clk_i clknet_leaf_59_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6006__A1 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8748_ _1048_ clknet_leaf_90_clk_i memory\[7\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7626__S _3806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8679_ _0979_ clknet_leaf_108_clk_i memory\[5\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3918__I1 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7361__S _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6493__A1 _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4985__S _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7293__I0 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6245__A1 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6705__S _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4225__S _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_51_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3909__I1 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3863__I net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5056__S _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ _1256_ memory\[18\]\[8\] _1376_ _1385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4582__I1 _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4291_ _1346_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6030_ _2629_ _2631_ _2495_ _2632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_60_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6484__A1 _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input5_I address_i[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7070__I _3505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6236__A1 _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7981_ _0281_ clknet_leaf_53_clk_i memory\[21\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_68_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6932_ _3443_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6863_ memory\[14\]\[9\] _1189_ _3397_ _3407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5814_ _1915_ _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7587__I1 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8602_ _0902_ clknet_leaf_208_clk_i memory\[4\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6794_ _3370_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5745_ _2163_ _2352_ _2029_ _2353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3974__S _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7446__S _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8533_ _0833_ clknet_leaf_200_clk_i memory\[8\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8464_ _0764_ clknet_leaf_60_clk_i memory\[31\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5676_ _1857_ _2281_ _2283_ _2284_ _2285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7415_ _1123_ memory\[0\]\[12\] _3697_ _3700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_79_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5474__B _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4627_ _1528_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_20_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8395_ _0695_ clknet_leaf_110_clk_i memory\[16\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6711__A2 _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7346_ _3663_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_92_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4558_ _1491_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7277_ _1121_ memory\[3\]\[11\] _3625_ _3627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4489_ _1454_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5921__C _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _1058_ _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6475__A1 _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6159_ _2753_ _2756_ _2757_ _2758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7275__I0 _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6227__B2 _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4109__I _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3948__I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_15_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6260__S _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6702__A2 _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput40 net40 data_o[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_102_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput51 net51 data_o[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput62 net62 data_o[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6466__A1 _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7266__I0 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6218__A1 _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5441__A2 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6662__C _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7569__I1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3860_ _1065_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_63_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7266__S _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4252__I0 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_119_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5530_ _1997_ _2139_ _2141_ _2142_ _2143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5461_ _1866_ _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4689__I _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7200_ _1112_ memory\[8\]\[7\] _3578_ _3586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4412_ _1412_ _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8180_ _0480_ clknet_leaf_35_clk_i memory\[27\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5392_ _2005_ _2007_ memory\[5\]\[1\] _2008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4555__I1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7131_ _3549_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4343_ _1375_ _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7062_ memory\[31\]\[6\] _1183_ _3506_ _3513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5741__C _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4274_ _1242_ memory\[17\]\[1\] _1336_ _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6013_ _2337_ _2526_ memory\[25\]\[15\] _2615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5313__I _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6209__A1 _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7964_ _0264_ clknet_leaf_40_clk_i memory\[20\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6915_ _1100_ memory\[16\]\[1\] _3433_ _3435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7895_ _0195_ clknet_leaf_29_clk_i memory\[18\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_25_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6846_ _3398_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4243__I0 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6777_ _1093_ memory\[9\]\[0\] _3361_ _3362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_135_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5916__C _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8516_ _0816_ clknet_leaf_118_clk_i memory\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3989_ memory\[19\]\[27\] _1154_ _1140_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5728_ _1862_ memory\[27\]\[9\] _2335_ _1867_ _2336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7176__S _3564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_189_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5659_ _2267_ memory\[1\]\[7\] _2268_ _2043_ _2269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8447_ _0747_ clknet_leaf_172_clk_i memory\[13\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_107_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4546__I1 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8378_ _0678_ clknet_leaf_216_clk_i memory\[14\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7329_ _3654_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5424__S _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5651__C _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7248__I0 _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6763__B _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_116_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3879__S _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5379__B _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6620__A1 _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4503__S _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4785__I1 _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_125_Left_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6687__A1 _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7487__I0 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6439__A1 _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_134_Left_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6611__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6392__C _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5965__A3 _2567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4961_ _1707_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4473__I0 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7680_ _1116_ memory\[7\]\[9\] _3837_ _3840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6700_ memory\[20\]\[30\] memory\[21\]\[30\] _1869_ _3287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4892_ _1089_ memory\[25\]\[30\] _1637_ _1671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3912_ memory\[19\]\[2\] _1102_ _1098_ _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7411__I0 _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4225__I0 _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6631_ memory\[8\]\[28\] memory\[9\]\[28\] _1992_ _3220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4413__S _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8301_ _0601_ clknet_leaf_58_clk_i net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6562_ _2846_ _3131_ _3151_ _3152_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_42_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4776__I1 _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_190_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6493_ _2674_ memory\[18\]\[25\] _3085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_15_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5308__I _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5513_ memory\[15\]\[4\] _1922_ _2125_ _1925_ _2126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_30_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8232_ _0532_ clknet_leaf_112_clk_i memory\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4528__I1 _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5444_ _1957_ memory\[26\]\[3\] _2058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8163_ _0463_ clknet_leaf_164_clk_i memory\[27\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5375_ _1987_ memory\[1\]\[1\] _1989_ _1990_ _1991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7114_ memory\[31\]\[31\] _1235_ _3505_ _3540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8094_ _0394_ clknet_leaf_19_clk_i memory\[24\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4326_ _1080_ memory\[17\]\[26\] _1358_ _1365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4257_ _1328_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7045_ memory\[13\]\[31\] _1235_ _3468_ _3503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_2_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4188_ _1084_ memory\[15\]\[28\] _1280_ _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_87_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7947_ _0247_ clknet_leaf_43_clk_i memory\[20\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7878_ _0178_ clknet_leaf_143_clk_i memory\[18\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7402__I0 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6829_ _1150_ memory\[9\]\[25\] _3383_ _3389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4216__I0 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5419__S _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7634__S _3806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4519__I1 _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6669__B2 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5662__B _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6758__B _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_129_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4455__I0 _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4233__S _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5556__C _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5580__A1 _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5572__B _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5332__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5064__S _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5291__C _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5160_ _1813_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5091_ _1082_ memory\[28\]\[27\] _1769_ _1777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4111_ _1239_ _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4042_ memory\[12\]\[10\] _1191_ _1192_ _1193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_137_clk_i_I clknet_4_9_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4694__I0 _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4408__S _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5993_ memory\[8\]\[14\] memory\[9\]\[14\] _2314_ _2596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4446__I0 _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5399__A1 _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7801_ _0101_ clknet_leaf_220_clk_i memory\[15\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6060__A2 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7732_ _0032_ clknet_leaf_28_clk_i memory\[19\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4944_ _1072_ memory\[26\]\[22\] _1696_ _1699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4875_ _1662_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7663_ _1100_ memory\[7\]\[1\] _1087_ _3831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4143__S _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7594_ _3794_ _3795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5466__C _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6614_ _3200_ _3202_ _1889_ _3203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5571__A1 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6545_ _2828_ memory\[10\]\[26\] _3136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7454__S _3685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8215_ _0515_ clknet_leaf_23_clk_i memory\[28\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6476_ _3053_ _3058_ _3063_ _3068_ _2894_ _3069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__7253__I _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5427_ _1988_ memory\[0\]\[2\] _2042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_100_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8146_ _0446_ clknet_leaf_43_clk_i memory\[26\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5358_ _1909_ _1973_ _1913_ _1974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8077_ _0377_ clknet_leaf_56_clk_i memory\[24\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4309_ _1277_ memory\[17\]\[18\] _1347_ _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5289_ _1905_ memory\[18\]\[0\] _1906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5626__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7028_ _3494_ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4318__S _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4988__I1 _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5149__S _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4988__S _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3892__S _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7364__S _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6488__B _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5314__A1 _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7539__S _3759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5567__B _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6670__C _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4979__I1 _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3866__I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ _1545_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4898__S _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_63_clk_i_I clknet_4_7_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4591_ _1508_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _2779_ _2925_ _2643_ _2926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6261_ _2754_ _2857_ _2666_ _2858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _2562_ memory\[6\]\[18\] _2791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8000_ _0300_ clknet_leaf_132_clk_i memory\[21\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5212_ _1818_ _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5143_ _1804_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5522__S _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5074_ _1056_ memory\[28\]\[19\] _1758_ _1768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4025_ net33 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_84_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7081__I1 _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3977__S _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4419__I0 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5976_ _2576_ _2578_ _2291_ _2579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4927_ _1269_ memory\[26\]\[14\] _1685_ _1690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5792__A1 _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7715_ _0015_ clknet_leaf_138_clk_i memory\[19\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8695_ _0995_ clknet_leaf_209_clk_i memory\[5\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4858_ _1653_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7646_ _3822_ _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4789_ memory\[24\]\[13\] _1198_ _1613_ _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4601__S _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7577_ memory\[5\]\[24\] net22 _3781_ _3786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6528_ memory\[30\]\[26\] memory\[31\]\[26\] _1923_ _3119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6459_ memory\[15\]\[24\] _2823_ _3051_ _2773_ _3052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__6895__I1 _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5940__B _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3858__A1 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8129_ _0429_ clknet_leaf_165_clk_i memory\[26\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6528__S _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4048__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7359__S _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5083__I0 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5783__A1 _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4830__I0 _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5535__A1 _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7094__S _3528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4511__S _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5838__A2 _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5830_ _2332_ _2431_ _2434_ _2435_ _2436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__6173__S _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5074__I0 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5761_ _2267_ memory\[1\]\[9\] _2368_ _2043_ _2369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_91_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5297__B _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ _1574_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8480_ _0780_ clknet_leaf_180_clk_i memory\[31\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7500_ _1139_ memory\[10\]\[20\] _3744_ _3745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6901__S _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5692_ _2163_ _2300_ _2029_ _2301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7431_ _3685_ _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_126_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4643_ memory\[22\]\[11\] _1194_ _1535_ _1537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5517__S _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4574_ memory\[21\]\[11\] _1194_ _1498_ _1500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4421__S _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7362_ _3671_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7293_ _1137_ memory\[3\]\[19\] _3625_ _3635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6313_ memory\[20\]\[21\] memory\[21\]\[21\] _2812_ _2909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5829__A2 _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6244_ _2472_ _2473_ memory\[5\]\[19\] _2842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_0_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4888__I0 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6175_ memory\[15\]\[18\] _2357_ _2772_ _2773_ _2774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5126_ _1263_ memory\[2\]\[11\] _1794_ _1796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5057_ _1759_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4008_ net38 _1168_ _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6591__B _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7054__I1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5959_ _2562_ memory\[6\]\[13\] _2563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8747_ _1047_ clknet_leaf_90_clk_i memory\[7\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8678_ _0978_ clknet_leaf_114_clk_i memory\[5\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_97_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7629_ _3813_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6868__I1 _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6485__C _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_11_clk_i_I clknet_4_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7089__S _3517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5056__I0 _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4008__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__I1 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5756__A1 _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__A1 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4241__S _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7552__S _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4040__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6859__I1 _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4290_ _1258_ memory\[17\]\[9\] _1336_ _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5072__S _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_173_clk_i clknet_4_8_0_clk_i clknet_leaf_173_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7980_ _0280_ clknet_leaf_52_clk_i memory\[21\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5800__S _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6931_ _1116_ memory\[16\]\[9\] _3433_ _3443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_188_clk_i clknet_4_3_0_clk_i clknet_leaf_188_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5047__I0 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6862_ _3406_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5813_ _2418_ _2419_ _2136_ _2420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_92_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8601_ _0901_ clknet_leaf_209_clk_i memory\[4\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6795__I0 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6793_ _1114_ memory\[9\]\[8\] _3361_ _3370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_111_clk_i clknet_4_15_0_clk_i clknet_leaf_111_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8532_ _0832_ clknet_leaf_80_clk_i memory\[8\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6631__S _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5744_ memory\[16\]\[9\] memory\[17\]\[9\] _2164_ _2352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8463_ _0763_ clknet_leaf_59_clk_i memory\[31\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7526__I _3758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5675_ _1871_ _2060_ memory\[25\]\[8\] _2284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_7414_ _3699_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8394_ _0694_ clknet_leaf_87_clk_i memory\[16\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_126_clk_i clknet_4_14_0_clk_i clknet_leaf_126_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_79_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4626_ memory\[22\]\[3\] _1177_ _1524_ _1528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_130_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7345_ _1121_ memory\[4\]\[11\] _3661_ _3663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_79_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4557_ memory\[21\]\[3\] _1177_ _1487_ _1491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7462__S _3722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7276_ _3626_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4488_ memory\[20\]\[3\] _1177_ _1450_ _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6227_ memory\[15\]\[19\] _2823_ _2824_ _2773_ _2825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_0_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6158_ _1889_ _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6227__A2 _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5109_ _1246_ memory\[2\]\[3\] _1783_ _1787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6806__S _3372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6089_ _2318_ memory\[0\]\[16\] _2690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_leaf_185_clk_i_I clknet_4_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5986__B2 _2588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4326__S _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7027__I1 _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7637__S _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4410__A1 _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5157__S _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4996__S _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6163__B2 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5210__I0 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7372__S _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput41 net41 data_o[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_leaf_90_clk_i clknet_4_13_0_clk_i clknet_leaf_90_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xoutput52 net52 data_o[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__6496__B _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput63 net63 data_o[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_47_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7018__I1 _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6777__I0 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_43_clk_i clknet_4_4_0_clk_i clknet_leaf_43_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6154__A1 _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5460_ _1905_ memory\[18\]\[3\] _2074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_54_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _1298_ _1411_ _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_41_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5901__A1 _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5391_ _2006_ _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_10_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_58_clk_i clknet_4_7_0_clk_i clknet_leaf_58_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7130_ memory\[11\]\[6\] _1183_ _3542_ _3549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4342_ _1095_ _1374_ _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7061_ _3512_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4273_ _1337_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6012_ _2382_ memory\[27\]\[15\] _2613_ _2384_ _2614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_74_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

