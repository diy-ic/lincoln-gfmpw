magic
tech gf180mcuD
magscale 1 10
timestamp 1701880005
<< obsm1 >>
rect 1344 3076 109984 111746
<< metal2 >>
rect 32928 114181 33040 114981
rect 33600 114181 33712 114981
rect 34272 114181 34384 114981
rect 36960 114181 37072 114981
rect 37632 114181 37744 114981
rect 38304 114181 38416 114981
rect 38976 114181 39088 114981
rect 46368 114181 46480 114981
rect 47040 114181 47152 114981
rect 47712 114181 47824 114981
rect 48384 114181 48496 114981
rect 50400 114181 50512 114981
rect 52416 114181 52528 114981
rect 55776 114181 55888 114981
rect 61152 114181 61264 114981
rect 63840 114181 63952 114981
rect 64512 114181 64624 114981
rect 68544 114181 68656 114981
rect 22176 0 22288 800
rect 32256 0 32368 800
rect 33600 0 33712 800
rect 34944 0 35056 800
rect 35616 0 35728 800
rect 47040 0 47152 800
rect 47712 0 47824 800
rect 53760 0 53872 800
rect 55104 0 55216 800
rect 61152 0 61264 800
rect 63168 0 63280 800
rect 64512 0 64624 800
rect 69888 0 70000 800
<< obsm2 >>
rect 1708 114121 32868 114181
rect 33100 114121 33540 114181
rect 33772 114121 34212 114181
rect 34444 114121 36900 114181
rect 37132 114121 37572 114181
rect 37804 114121 38244 114181
rect 38476 114121 38916 114181
rect 39148 114121 46308 114181
rect 46540 114121 46980 114181
rect 47212 114121 47652 114181
rect 47884 114121 48324 114181
rect 48556 114121 50340 114181
rect 50572 114121 52356 114181
rect 52588 114121 55716 114181
rect 55948 114121 61092 114181
rect 61324 114121 63780 114181
rect 64012 114121 64452 114181
rect 64684 114121 68484 114181
rect 68716 114121 110740 114181
rect 1708 860 110740 114121
rect 1708 700 22116 860
rect 22348 700 32196 860
rect 32428 700 33540 860
rect 33772 700 34884 860
rect 35116 700 35556 860
rect 35788 700 46980 860
rect 47212 700 47652 860
rect 47884 700 53700 860
rect 53932 700 55044 860
rect 55276 700 61092 860
rect 61324 700 63108 860
rect 63340 700 64452 860
rect 64684 700 69828 860
rect 70060 700 110740 860
<< metal3 >>
rect 0 109536 800 109648
rect 110597 81984 111397 82096
rect 0 79296 800 79408
rect 110597 79296 111397 79408
rect 110597 78624 111397 78736
rect 110597 71232 111397 71344
rect 0 70560 800 70672
rect 110597 70560 111397 70672
rect 110597 69216 111397 69328
rect 0 68544 800 68656
rect 110597 67200 111397 67312
rect 110597 66528 111397 66640
rect 110597 64512 111397 64624
rect 110597 63168 111397 63280
rect 0 62496 800 62608
rect 110597 62496 111397 62608
rect 0 59808 800 59920
rect 0 58464 800 58576
rect 110597 57792 111397 57904
rect 0 57120 800 57232
rect 110597 57120 111397 57232
rect 110597 53088 111397 53200
rect 110597 52416 111397 52528
rect 110597 51744 111397 51856
rect 110597 48384 111397 48496
rect 110597 43008 111397 43120
rect 110597 42336 111397 42448
rect 110597 41664 111397 41776
rect 0 38976 800 39088
rect 0 38304 800 38416
rect 0 37632 800 37744
rect 0 36960 800 37072
rect 0 36288 800 36400
rect 0 34944 800 35056
rect 0 34272 800 34384
rect 0 33600 800 33712
rect 0 31584 800 31696
rect 0 28896 800 29008
rect 0 25536 800 25648
rect 0 22848 800 22960
<< obsm3 >>
rect 800 109708 110740 112532
rect 860 109476 110740 109708
rect 800 82156 110740 109476
rect 800 81924 110537 82156
rect 800 79468 110740 81924
rect 860 79236 110537 79468
rect 800 78796 110740 79236
rect 800 78564 110537 78796
rect 800 71404 110740 78564
rect 800 71172 110537 71404
rect 800 70732 110740 71172
rect 860 70500 110537 70732
rect 800 69388 110740 70500
rect 800 69156 110537 69388
rect 800 68716 110740 69156
rect 860 68484 110740 68716
rect 800 67372 110740 68484
rect 800 67140 110537 67372
rect 800 66700 110740 67140
rect 800 66468 110537 66700
rect 800 64684 110740 66468
rect 800 64452 110537 64684
rect 800 63340 110740 64452
rect 800 63108 110537 63340
rect 800 62668 110740 63108
rect 860 62436 110537 62668
rect 800 59980 110740 62436
rect 860 59748 110740 59980
rect 800 58636 110740 59748
rect 860 58404 110740 58636
rect 800 57964 110740 58404
rect 800 57732 110537 57964
rect 800 57292 110740 57732
rect 860 57060 110537 57292
rect 800 53260 110740 57060
rect 800 53028 110537 53260
rect 800 52588 110740 53028
rect 800 52356 110537 52588
rect 800 51916 110740 52356
rect 800 51684 110537 51916
rect 800 48556 110740 51684
rect 800 48324 110537 48556
rect 800 43180 110740 48324
rect 800 42948 110537 43180
rect 800 42508 110740 42948
rect 800 42276 110537 42508
rect 800 41836 110740 42276
rect 800 41604 110537 41836
rect 800 39148 110740 41604
rect 860 38916 110740 39148
rect 800 38476 110740 38916
rect 860 38244 110740 38476
rect 800 37804 110740 38244
rect 860 37572 110740 37804
rect 800 37132 110740 37572
rect 860 36900 110740 37132
rect 800 36460 110740 36900
rect 860 36228 110740 36460
rect 800 35116 110740 36228
rect 860 34884 110740 35116
rect 800 34444 110740 34884
rect 860 34212 110740 34444
rect 800 33772 110740 34212
rect 860 33540 110740 33772
rect 800 31756 110740 33540
rect 860 31524 110740 31756
rect 800 29068 110740 31524
rect 860 28836 110740 29068
rect 800 25708 110740 28836
rect 860 25476 110740 25708
rect 800 23020 110740 25476
rect 860 22788 110740 23020
rect 800 3108 110740 22788
<< metal4 >>
rect 4448 3076 4768 111388
rect 19808 3076 20128 111388
rect 35168 3076 35488 111388
rect 50528 3076 50848 111388
rect 65888 3076 66208 111388
rect 81248 3076 81568 111388
rect 96608 3076 96928 111388
<< obsm4 >>
rect 1932 3266 4388 110974
rect 4828 3266 19748 110974
rect 20188 3266 35108 110974
rect 35548 3266 50468 110974
rect 50908 3266 65828 110974
rect 66268 3266 81188 110974
rect 81628 3266 96548 110974
rect 96988 3266 109508 110974
<< labels >>
rlabel metal3 s 0 62496 800 62608 6 address_i[0]
port 1 nsew signal input
rlabel metal3 s 0 58464 800 58576 6 address_i[1]
port 2 nsew signal input
rlabel metal3 s 0 57120 800 57232 6 address_i[2]
port 3 nsew signal input
rlabel metal3 s 110597 57120 111397 57232 6 address_i[3]
port 4 nsew signal input
rlabel metal2 s 61152 0 61264 800 6 address_i[4]
port 5 nsew signal input
rlabel metal3 s 0 109536 800 109648 6 clk_i
port 6 nsew signal input
rlabel metal3 s 110597 51744 111397 51856 6 data_i[0]
port 7 nsew signal input
rlabel metal2 s 63840 114181 63952 114981 6 data_i[10]
port 8 nsew signal input
rlabel metal2 s 64512 114181 64624 114981 6 data_i[11]
port 9 nsew signal input
rlabel metal2 s 61152 114181 61264 114981 6 data_i[12]
port 10 nsew signal input
rlabel metal2 s 55776 114181 55888 114981 6 data_i[13]
port 11 nsew signal input
rlabel metal2 s 52416 114181 52528 114981 6 data_i[14]
port 12 nsew signal input
rlabel metal2 s 47040 114181 47152 114981 6 data_i[15]
port 13 nsew signal input
rlabel metal2 s 47712 114181 47824 114981 6 data_i[16]
port 14 nsew signal input
rlabel metal2 s 46368 114181 46480 114981 6 data_i[17]
port 15 nsew signal input
rlabel metal2 s 50400 114181 50512 114981 6 data_i[18]
port 16 nsew signal input
rlabel metal2 s 48384 114181 48496 114981 6 data_i[19]
port 17 nsew signal input
rlabel metal3 s 110597 52416 111397 52528 6 data_i[1]
port 18 nsew signal input
rlabel metal2 s 47712 0 47824 800 6 data_i[20]
port 19 nsew signal input
rlabel metal2 s 35616 0 35728 800 6 data_i[21]
port 20 nsew signal input
rlabel metal2 s 32256 0 32368 800 6 data_i[22]
port 21 nsew signal input
rlabel metal3 s 0 28896 800 29008 6 data_i[23]
port 22 nsew signal input
rlabel metal3 s 0 25536 800 25648 6 data_i[24]
port 23 nsew signal input
rlabel metal2 s 22176 0 22288 800 6 data_i[25]
port 24 nsew signal input
rlabel metal3 s 0 22848 800 22960 6 data_i[26]
port 25 nsew signal input
rlabel metal3 s 0 31584 800 31696 6 data_i[27]
port 26 nsew signal input
rlabel metal2 s 47040 0 47152 800 6 data_i[28]
port 27 nsew signal input
rlabel metal2 s 53760 0 53872 800 6 data_i[29]
port 28 nsew signal input
rlabel metal3 s 110597 53088 111397 53200 6 data_i[2]
port 29 nsew signal input
rlabel metal2 s 55104 0 55216 800 6 data_i[30]
port 30 nsew signal input
rlabel metal2 s 63168 0 63280 800 6 data_i[31]
port 31 nsew signal input
rlabel metal3 s 110597 57792 111397 57904 6 data_i[3]
port 32 nsew signal input
rlabel metal3 s 110597 62496 111397 62608 6 data_i[4]
port 33 nsew signal input
rlabel metal3 s 110597 71232 111397 71344 6 data_i[5]
port 34 nsew signal input
rlabel metal3 s 110597 78624 111397 78736 6 data_i[6]
port 35 nsew signal input
rlabel metal3 s 110597 81984 111397 82096 6 data_i[7]
port 36 nsew signal input
rlabel metal3 s 110597 79296 111397 79408 6 data_i[8]
port 37 nsew signal input
rlabel metal2 s 68544 114181 68656 114981 6 data_i[9]
port 38 nsew signal input
rlabel metal3 s 110597 42336 111397 42448 6 data_o[0]
port 39 nsew signal output
rlabel metal2 s 38304 114181 38416 114981 6 data_o[10]
port 40 nsew signal output
rlabel metal2 s 37632 114181 37744 114981 6 data_o[11]
port 41 nsew signal output
rlabel metal2 s 36960 114181 37072 114981 6 data_o[12]
port 42 nsew signal output
rlabel metal2 s 34272 114181 34384 114981 6 data_o[13]
port 43 nsew signal output
rlabel metal2 s 33600 114181 33712 114981 6 data_o[14]
port 44 nsew signal output
rlabel metal2 s 32928 114181 33040 114981 6 data_o[15]
port 45 nsew signal output
rlabel metal2 s 38976 114181 39088 114981 6 data_o[16]
port 46 nsew signal output
rlabel metal3 s 0 79296 800 79408 6 data_o[17]
port 47 nsew signal output
rlabel metal3 s 0 70560 800 70672 6 data_o[18]
port 48 nsew signal output
rlabel metal3 s 0 68544 800 68656 6 data_o[19]
port 49 nsew signal output
rlabel metal3 s 110597 43008 111397 43120 6 data_o[1]
port 50 nsew signal output
rlabel metal2 s 34944 0 35056 800 6 data_o[20]
port 51 nsew signal output
rlabel metal3 s 0 36288 800 36400 6 data_o[21]
port 52 nsew signal output
rlabel metal2 s 33600 0 33712 800 6 data_o[22]
port 53 nsew signal output
rlabel metal3 s 0 34944 800 35056 6 data_o[23]
port 54 nsew signal output
rlabel metal3 s 0 34272 800 34384 6 data_o[24]
port 55 nsew signal output
rlabel metal3 s 0 37632 800 37744 6 data_o[25]
port 56 nsew signal output
rlabel metal3 s 0 38976 800 39088 6 data_o[26]
port 57 nsew signal output
rlabel metal3 s 0 33600 800 33712 6 data_o[27]
port 58 nsew signal output
rlabel metal3 s 0 36960 800 37072 6 data_o[28]
port 59 nsew signal output
rlabel metal3 s 0 38304 800 38416 6 data_o[29]
port 60 nsew signal output
rlabel metal3 s 110597 41664 111397 41776 6 data_o[2]
port 61 nsew signal output
rlabel metal2 s 64512 0 64624 800 6 data_o[30]
port 62 nsew signal output
rlabel metal2 s 69888 0 70000 800 6 data_o[31]
port 63 nsew signal output
rlabel metal3 s 110597 48384 111397 48496 6 data_o[3]
port 64 nsew signal output
rlabel metal3 s 110597 63168 111397 63280 6 data_o[4]
port 65 nsew signal output
rlabel metal3 s 110597 64512 111397 64624 6 data_o[5]
port 66 nsew signal output
rlabel metal3 s 110597 67200 111397 67312 6 data_o[6]
port 67 nsew signal output
rlabel metal3 s 110597 66528 111397 66640 6 data_o[7]
port 68 nsew signal output
rlabel metal3 s 110597 69216 111397 69328 6 data_o[8]
port 69 nsew signal output
rlabel metal3 s 110597 70560 111397 70672 6 data_o[9]
port 70 nsew signal output
rlabel metal4 s 4448 3076 4768 111388 6 vdd
port 71 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 111388 6 vdd
port 71 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 111388 6 vdd
port 71 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 111388 6 vdd
port 71 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 111388 6 vss
port 72 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 111388 6 vss
port 72 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 111388 6 vss
port 72 nsew ground bidirectional
rlabel metal3 s 0 59808 800 59920 6 we_i
port 73 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 111397 114981
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10683626
string GDS_FILE /home/kris/repos/diy-ic/lincoln-gfmpw/openlane/ram_block/runs/23_12_06_16_20/results/signoff/ram.magic.gds
string GDS_START 260750
<< end >>

