magic
tech gf180mcuD
magscale 1 5
timestamp 1702002516
<< obsm1 >>
rect 672 855 79296 78430
<< metal2 >>
rect 7616 0 7672 400
rect 7952 0 8008 400
rect 8288 0 8344 400
rect 8624 0 8680 400
rect 8960 0 9016 400
rect 9296 0 9352 400
rect 9632 0 9688 400
rect 9968 0 10024 400
rect 10304 0 10360 400
rect 10640 0 10696 400
rect 10976 0 11032 400
rect 11312 0 11368 400
rect 11648 0 11704 400
rect 11984 0 12040 400
rect 12320 0 12376 400
rect 12656 0 12712 400
rect 12992 0 13048 400
rect 13328 0 13384 400
rect 13664 0 13720 400
rect 14000 0 14056 400
rect 14336 0 14392 400
rect 14672 0 14728 400
rect 15008 0 15064 400
rect 15344 0 15400 400
rect 15680 0 15736 400
rect 16016 0 16072 400
rect 16352 0 16408 400
rect 16688 0 16744 400
rect 17024 0 17080 400
rect 17360 0 17416 400
rect 17696 0 17752 400
rect 18032 0 18088 400
rect 18368 0 18424 400
rect 18704 0 18760 400
rect 19040 0 19096 400
rect 19376 0 19432 400
rect 19712 0 19768 400
rect 20048 0 20104 400
rect 20384 0 20440 400
rect 20720 0 20776 400
rect 21056 0 21112 400
rect 21392 0 21448 400
rect 21728 0 21784 400
rect 22064 0 22120 400
rect 22400 0 22456 400
rect 22736 0 22792 400
rect 23072 0 23128 400
rect 23408 0 23464 400
rect 23744 0 23800 400
rect 24080 0 24136 400
rect 24416 0 24472 400
rect 24752 0 24808 400
rect 25088 0 25144 400
rect 25424 0 25480 400
rect 25760 0 25816 400
rect 26096 0 26152 400
rect 26432 0 26488 400
rect 26768 0 26824 400
rect 27104 0 27160 400
rect 27440 0 27496 400
rect 27776 0 27832 400
rect 28112 0 28168 400
rect 28448 0 28504 400
rect 28784 0 28840 400
rect 29120 0 29176 400
rect 29456 0 29512 400
rect 29792 0 29848 400
rect 30128 0 30184 400
rect 30464 0 30520 400
rect 30800 0 30856 400
rect 31136 0 31192 400
rect 31472 0 31528 400
rect 31808 0 31864 400
rect 32144 0 32200 400
rect 32480 0 32536 400
rect 32816 0 32872 400
rect 33152 0 33208 400
rect 33488 0 33544 400
rect 33824 0 33880 400
rect 34160 0 34216 400
rect 34496 0 34552 400
rect 34832 0 34888 400
rect 35168 0 35224 400
rect 35504 0 35560 400
rect 35840 0 35896 400
rect 36176 0 36232 400
rect 36512 0 36568 400
rect 36848 0 36904 400
rect 37184 0 37240 400
rect 37520 0 37576 400
rect 37856 0 37912 400
rect 38192 0 38248 400
rect 38528 0 38584 400
rect 38864 0 38920 400
rect 39200 0 39256 400
rect 39536 0 39592 400
rect 39872 0 39928 400
rect 40208 0 40264 400
rect 40544 0 40600 400
rect 40880 0 40936 400
rect 41216 0 41272 400
rect 41552 0 41608 400
rect 41888 0 41944 400
rect 42224 0 42280 400
rect 42560 0 42616 400
rect 42896 0 42952 400
rect 43232 0 43288 400
rect 43568 0 43624 400
rect 43904 0 43960 400
rect 44240 0 44296 400
rect 44576 0 44632 400
rect 44912 0 44968 400
rect 45248 0 45304 400
rect 45584 0 45640 400
rect 45920 0 45976 400
rect 46256 0 46312 400
rect 46592 0 46648 400
rect 46928 0 46984 400
rect 47264 0 47320 400
rect 47600 0 47656 400
rect 47936 0 47992 400
rect 48272 0 48328 400
rect 48608 0 48664 400
rect 48944 0 49000 400
rect 49280 0 49336 400
rect 49616 0 49672 400
rect 49952 0 50008 400
rect 50288 0 50344 400
rect 50624 0 50680 400
rect 50960 0 51016 400
rect 51296 0 51352 400
rect 51632 0 51688 400
rect 51968 0 52024 400
rect 52304 0 52360 400
rect 52640 0 52696 400
rect 52976 0 53032 400
rect 53312 0 53368 400
rect 53648 0 53704 400
rect 53984 0 54040 400
rect 54320 0 54376 400
rect 54656 0 54712 400
rect 54992 0 55048 400
rect 55328 0 55384 400
rect 55664 0 55720 400
rect 56000 0 56056 400
rect 56336 0 56392 400
rect 56672 0 56728 400
rect 57008 0 57064 400
rect 57344 0 57400 400
rect 57680 0 57736 400
rect 58016 0 58072 400
rect 58352 0 58408 400
rect 58688 0 58744 400
rect 59024 0 59080 400
rect 59360 0 59416 400
rect 59696 0 59752 400
rect 60032 0 60088 400
rect 60368 0 60424 400
rect 60704 0 60760 400
rect 61040 0 61096 400
rect 61376 0 61432 400
rect 61712 0 61768 400
rect 62048 0 62104 400
rect 62384 0 62440 400
rect 62720 0 62776 400
rect 63056 0 63112 400
rect 63392 0 63448 400
rect 63728 0 63784 400
rect 64064 0 64120 400
rect 64400 0 64456 400
rect 64736 0 64792 400
rect 65072 0 65128 400
rect 65408 0 65464 400
rect 65744 0 65800 400
rect 66080 0 66136 400
rect 66416 0 66472 400
rect 66752 0 66808 400
rect 67088 0 67144 400
rect 67424 0 67480 400
rect 67760 0 67816 400
rect 68096 0 68152 400
rect 68432 0 68488 400
rect 68768 0 68824 400
rect 69104 0 69160 400
rect 69440 0 69496 400
rect 69776 0 69832 400
rect 70112 0 70168 400
rect 70448 0 70504 400
rect 70784 0 70840 400
rect 71120 0 71176 400
rect 71456 0 71512 400
rect 71792 0 71848 400
rect 72128 0 72184 400
<< obsm2 >>
rect 854 430 79282 78419
rect 854 400 7586 430
rect 7702 400 7922 430
rect 8038 400 8258 430
rect 8374 400 8594 430
rect 8710 400 8930 430
rect 9046 400 9266 430
rect 9382 400 9602 430
rect 9718 400 9938 430
rect 10054 400 10274 430
rect 10390 400 10610 430
rect 10726 400 10946 430
rect 11062 400 11282 430
rect 11398 400 11618 430
rect 11734 400 11954 430
rect 12070 400 12290 430
rect 12406 400 12626 430
rect 12742 400 12962 430
rect 13078 400 13298 430
rect 13414 400 13634 430
rect 13750 400 13970 430
rect 14086 400 14306 430
rect 14422 400 14642 430
rect 14758 400 14978 430
rect 15094 400 15314 430
rect 15430 400 15650 430
rect 15766 400 15986 430
rect 16102 400 16322 430
rect 16438 400 16658 430
rect 16774 400 16994 430
rect 17110 400 17330 430
rect 17446 400 17666 430
rect 17782 400 18002 430
rect 18118 400 18338 430
rect 18454 400 18674 430
rect 18790 400 19010 430
rect 19126 400 19346 430
rect 19462 400 19682 430
rect 19798 400 20018 430
rect 20134 400 20354 430
rect 20470 400 20690 430
rect 20806 400 21026 430
rect 21142 400 21362 430
rect 21478 400 21698 430
rect 21814 400 22034 430
rect 22150 400 22370 430
rect 22486 400 22706 430
rect 22822 400 23042 430
rect 23158 400 23378 430
rect 23494 400 23714 430
rect 23830 400 24050 430
rect 24166 400 24386 430
rect 24502 400 24722 430
rect 24838 400 25058 430
rect 25174 400 25394 430
rect 25510 400 25730 430
rect 25846 400 26066 430
rect 26182 400 26402 430
rect 26518 400 26738 430
rect 26854 400 27074 430
rect 27190 400 27410 430
rect 27526 400 27746 430
rect 27862 400 28082 430
rect 28198 400 28418 430
rect 28534 400 28754 430
rect 28870 400 29090 430
rect 29206 400 29426 430
rect 29542 400 29762 430
rect 29878 400 30098 430
rect 30214 400 30434 430
rect 30550 400 30770 430
rect 30886 400 31106 430
rect 31222 400 31442 430
rect 31558 400 31778 430
rect 31894 400 32114 430
rect 32230 400 32450 430
rect 32566 400 32786 430
rect 32902 400 33122 430
rect 33238 400 33458 430
rect 33574 400 33794 430
rect 33910 400 34130 430
rect 34246 400 34466 430
rect 34582 400 34802 430
rect 34918 400 35138 430
rect 35254 400 35474 430
rect 35590 400 35810 430
rect 35926 400 36146 430
rect 36262 400 36482 430
rect 36598 400 36818 430
rect 36934 400 37154 430
rect 37270 400 37490 430
rect 37606 400 37826 430
rect 37942 400 38162 430
rect 38278 400 38498 430
rect 38614 400 38834 430
rect 38950 400 39170 430
rect 39286 400 39506 430
rect 39622 400 39842 430
rect 39958 400 40178 430
rect 40294 400 40514 430
rect 40630 400 40850 430
rect 40966 400 41186 430
rect 41302 400 41522 430
rect 41638 400 41858 430
rect 41974 400 42194 430
rect 42310 400 42530 430
rect 42646 400 42866 430
rect 42982 400 43202 430
rect 43318 400 43538 430
rect 43654 400 43874 430
rect 43990 400 44210 430
rect 44326 400 44546 430
rect 44662 400 44882 430
rect 44998 400 45218 430
rect 45334 400 45554 430
rect 45670 400 45890 430
rect 46006 400 46226 430
rect 46342 400 46562 430
rect 46678 400 46898 430
rect 47014 400 47234 430
rect 47350 400 47570 430
rect 47686 400 47906 430
rect 48022 400 48242 430
rect 48358 400 48578 430
rect 48694 400 48914 430
rect 49030 400 49250 430
rect 49366 400 49586 430
rect 49702 400 49922 430
rect 50038 400 50258 430
rect 50374 400 50594 430
rect 50710 400 50930 430
rect 51046 400 51266 430
rect 51382 400 51602 430
rect 51718 400 51938 430
rect 52054 400 52274 430
rect 52390 400 52610 430
rect 52726 400 52946 430
rect 53062 400 53282 430
rect 53398 400 53618 430
rect 53734 400 53954 430
rect 54070 400 54290 430
rect 54406 400 54626 430
rect 54742 400 54962 430
rect 55078 400 55298 430
rect 55414 400 55634 430
rect 55750 400 55970 430
rect 56086 400 56306 430
rect 56422 400 56642 430
rect 56758 400 56978 430
rect 57094 400 57314 430
rect 57430 400 57650 430
rect 57766 400 57986 430
rect 58102 400 58322 430
rect 58438 400 58658 430
rect 58774 400 58994 430
rect 59110 400 59330 430
rect 59446 400 59666 430
rect 59782 400 60002 430
rect 60118 400 60338 430
rect 60454 400 60674 430
rect 60790 400 61010 430
rect 61126 400 61346 430
rect 61462 400 61682 430
rect 61798 400 62018 430
rect 62134 400 62354 430
rect 62470 400 62690 430
rect 62806 400 63026 430
rect 63142 400 63362 430
rect 63478 400 63698 430
rect 63814 400 64034 430
rect 64150 400 64370 430
rect 64486 400 64706 430
rect 64822 400 65042 430
rect 65158 400 65378 430
rect 65494 400 65714 430
rect 65830 400 66050 430
rect 66166 400 66386 430
rect 66502 400 66722 430
rect 66838 400 67058 430
rect 67174 400 67394 430
rect 67510 400 67730 430
rect 67846 400 68066 430
rect 68182 400 68402 430
rect 68518 400 68738 430
rect 68854 400 69074 430
rect 69190 400 69410 430
rect 69526 400 69746 430
rect 69862 400 70082 430
rect 70198 400 70418 430
rect 70534 400 70754 430
rect 70870 400 71090 430
rect 71206 400 71426 430
rect 71542 400 71762 430
rect 71878 400 72098 430
rect 72214 400 79282 430
<< metal3 >>
rect 0 77280 400 77336
rect 79600 77280 80000 77336
rect 0 74032 400 74088
rect 79600 74032 80000 74088
rect 0 70784 400 70840
rect 79600 70784 80000 70840
rect 0 67536 400 67592
rect 79600 67536 80000 67592
rect 0 64288 400 64344
rect 79600 64288 80000 64344
rect 0 61040 400 61096
rect 79600 61040 80000 61096
rect 0 57792 400 57848
rect 79600 57792 80000 57848
rect 0 54544 400 54600
rect 79600 54544 80000 54600
rect 0 51296 400 51352
rect 79600 51296 80000 51352
rect 0 48048 400 48104
rect 79600 48048 80000 48104
rect 0 44800 400 44856
rect 79600 44800 80000 44856
rect 0 41552 400 41608
rect 79600 41552 80000 41608
rect 0 38304 400 38360
rect 79600 38304 80000 38360
rect 0 35056 400 35112
rect 79600 35056 80000 35112
rect 0 31808 400 31864
rect 79600 31808 80000 31864
rect 0 28560 400 28616
rect 79600 28560 80000 28616
rect 0 25312 400 25368
rect 79600 25312 80000 25368
rect 0 22064 400 22120
rect 79600 22064 80000 22120
rect 0 18816 400 18872
rect 79600 18816 80000 18872
rect 0 15568 400 15624
rect 79600 15568 80000 15624
rect 0 12320 400 12376
rect 79600 12320 80000 12376
rect 0 9072 400 9128
rect 79600 9072 80000 9128
rect 0 5824 400 5880
rect 79600 5824 80000 5880
rect 0 2576 400 2632
rect 79600 2576 80000 2632
<< obsm3 >>
rect 400 77366 79600 78414
rect 430 77250 79570 77366
rect 400 74118 79600 77250
rect 430 74002 79570 74118
rect 400 70870 79600 74002
rect 430 70754 79570 70870
rect 400 67622 79600 70754
rect 430 67506 79570 67622
rect 400 64374 79600 67506
rect 430 64258 79570 64374
rect 400 61126 79600 64258
rect 430 61010 79570 61126
rect 400 57878 79600 61010
rect 430 57762 79570 57878
rect 400 54630 79600 57762
rect 430 54514 79570 54630
rect 400 51382 79600 54514
rect 430 51266 79570 51382
rect 400 48134 79600 51266
rect 430 48018 79570 48134
rect 400 44886 79600 48018
rect 430 44770 79570 44886
rect 400 41638 79600 44770
rect 430 41522 79570 41638
rect 400 38390 79600 41522
rect 430 38274 79570 38390
rect 400 35142 79600 38274
rect 430 35026 79570 35142
rect 400 31894 79600 35026
rect 430 31778 79570 31894
rect 400 28646 79600 31778
rect 430 28530 79570 28646
rect 400 25398 79600 28530
rect 430 25282 79570 25398
rect 400 22150 79600 25282
rect 430 22034 79570 22150
rect 400 18902 79600 22034
rect 430 18786 79570 18902
rect 400 15654 79600 18786
rect 430 15538 79570 15654
rect 400 12406 79600 15538
rect 430 12290 79570 12406
rect 400 9158 79600 12290
rect 430 9042 79570 9158
rect 400 5910 79600 9042
rect 430 5794 79570 5910
rect 400 2662 79600 5794
rect 430 2546 79570 2662
rect 400 1470 79600 2546
<< metal4 >>
rect 2224 1538 2384 78430
rect 9904 1538 10064 78430
rect 17584 1538 17744 78430
rect 25264 1538 25424 78430
rect 32944 1538 33104 78430
rect 40624 1538 40784 78430
rect 48304 1538 48464 78430
rect 55984 1538 56144 78430
rect 63664 1538 63824 78430
rect 71344 1538 71504 78430
rect 79024 1538 79184 78430
<< obsm4 >>
rect 10486 2417 17554 59799
rect 17774 2417 25234 59799
rect 25454 2417 32914 59799
rect 33134 2417 40594 59799
rect 40814 2417 48274 59799
rect 48494 2417 55954 59799
rect 56174 2417 63634 59799
rect 63854 2417 66346 59799
<< labels >>
rlabel metal3 s 79600 2576 80000 2632 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 57792 400 57848 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 48048 400 48104 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 38304 400 38360 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 28560 400 28616 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 18816 400 18872 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 9072 400 9128 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 79600 12320 80000 12376 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 79600 22064 80000 22120 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 79600 31808 80000 31864 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 79600 41552 80000 41608 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 79600 51296 80000 51352 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 79600 61040 80000 61096 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 79600 70784 80000 70840 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 77280 400 77336 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 67536 400 67592 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 79600 9072 80000 9128 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 51296 400 51352 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 41552 400 41608 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 31808 400 31864 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 22064 400 22120 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 12320 400 12376 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 2576 400 2632 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 79600 18816 80000 18872 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 79600 28560 80000 28616 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 79600 38304 80000 38360 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 79600 48048 80000 48104 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 79600 57792 80000 57848 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 79600 67536 80000 67592 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 79600 77280 80000 77336 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 70784 400 70840 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 61040 400 61096 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 79600 5824 80000 5880 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 54544 400 54600 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 44800 400 44856 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 35056 400 35112 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 25312 400 25368 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 15568 400 15624 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 5824 400 5880 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 79600 15568 80000 15624 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 79600 25312 80000 25368 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 79600 35056 80000 35112 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 79600 44800 80000 44856 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 79600 54544 80000 54600 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 79600 64288 80000 64344 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 79600 74032 80000 74088 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 74032 400 74088 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 64288 400 64344 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 7952 0 8008 400 6 la_data_in[0]
port 49 nsew signal input
rlabel metal2 s 18032 0 18088 400 6 la_data_in[10]
port 50 nsew signal input
rlabel metal2 s 19040 0 19096 400 6 la_data_in[11]
port 51 nsew signal input
rlabel metal2 s 20048 0 20104 400 6 la_data_in[12]
port 52 nsew signal input
rlabel metal2 s 21056 0 21112 400 6 la_data_in[13]
port 53 nsew signal input
rlabel metal2 s 22064 0 22120 400 6 la_data_in[14]
port 54 nsew signal input
rlabel metal2 s 23072 0 23128 400 6 la_data_in[15]
port 55 nsew signal input
rlabel metal2 s 24080 0 24136 400 6 la_data_in[16]
port 56 nsew signal input
rlabel metal2 s 25088 0 25144 400 6 la_data_in[17]
port 57 nsew signal input
rlabel metal2 s 26096 0 26152 400 6 la_data_in[18]
port 58 nsew signal input
rlabel metal2 s 27104 0 27160 400 6 la_data_in[19]
port 59 nsew signal input
rlabel metal2 s 8960 0 9016 400 6 la_data_in[1]
port 60 nsew signal input
rlabel metal2 s 28112 0 28168 400 6 la_data_in[20]
port 61 nsew signal input
rlabel metal2 s 29120 0 29176 400 6 la_data_in[21]
port 62 nsew signal input
rlabel metal2 s 30128 0 30184 400 6 la_data_in[22]
port 63 nsew signal input
rlabel metal2 s 31136 0 31192 400 6 la_data_in[23]
port 64 nsew signal input
rlabel metal2 s 32144 0 32200 400 6 la_data_in[24]
port 65 nsew signal input
rlabel metal2 s 33152 0 33208 400 6 la_data_in[25]
port 66 nsew signal input
rlabel metal2 s 34160 0 34216 400 6 la_data_in[26]
port 67 nsew signal input
rlabel metal2 s 35168 0 35224 400 6 la_data_in[27]
port 68 nsew signal input
rlabel metal2 s 36176 0 36232 400 6 la_data_in[28]
port 69 nsew signal input
rlabel metal2 s 37184 0 37240 400 6 la_data_in[29]
port 70 nsew signal input
rlabel metal2 s 9968 0 10024 400 6 la_data_in[2]
port 71 nsew signal input
rlabel metal2 s 38192 0 38248 400 6 la_data_in[30]
port 72 nsew signal input
rlabel metal2 s 39200 0 39256 400 6 la_data_in[31]
port 73 nsew signal input
rlabel metal2 s 40208 0 40264 400 6 la_data_in[32]
port 74 nsew signal input
rlabel metal2 s 41216 0 41272 400 6 la_data_in[33]
port 75 nsew signal input
rlabel metal2 s 42224 0 42280 400 6 la_data_in[34]
port 76 nsew signal input
rlabel metal2 s 43232 0 43288 400 6 la_data_in[35]
port 77 nsew signal input
rlabel metal2 s 44240 0 44296 400 6 la_data_in[36]
port 78 nsew signal input
rlabel metal2 s 45248 0 45304 400 6 la_data_in[37]
port 79 nsew signal input
rlabel metal2 s 46256 0 46312 400 6 la_data_in[38]
port 80 nsew signal input
rlabel metal2 s 47264 0 47320 400 6 la_data_in[39]
port 81 nsew signal input
rlabel metal2 s 10976 0 11032 400 6 la_data_in[3]
port 82 nsew signal input
rlabel metal2 s 48272 0 48328 400 6 la_data_in[40]
port 83 nsew signal input
rlabel metal2 s 49280 0 49336 400 6 la_data_in[41]
port 84 nsew signal input
rlabel metal2 s 50288 0 50344 400 6 la_data_in[42]
port 85 nsew signal input
rlabel metal2 s 51296 0 51352 400 6 la_data_in[43]
port 86 nsew signal input
rlabel metal2 s 52304 0 52360 400 6 la_data_in[44]
port 87 nsew signal input
rlabel metal2 s 53312 0 53368 400 6 la_data_in[45]
port 88 nsew signal input
rlabel metal2 s 54320 0 54376 400 6 la_data_in[46]
port 89 nsew signal input
rlabel metal2 s 55328 0 55384 400 6 la_data_in[47]
port 90 nsew signal input
rlabel metal2 s 56336 0 56392 400 6 la_data_in[48]
port 91 nsew signal input
rlabel metal2 s 57344 0 57400 400 6 la_data_in[49]
port 92 nsew signal input
rlabel metal2 s 11984 0 12040 400 6 la_data_in[4]
port 93 nsew signal input
rlabel metal2 s 58352 0 58408 400 6 la_data_in[50]
port 94 nsew signal input
rlabel metal2 s 59360 0 59416 400 6 la_data_in[51]
port 95 nsew signal input
rlabel metal2 s 60368 0 60424 400 6 la_data_in[52]
port 96 nsew signal input
rlabel metal2 s 61376 0 61432 400 6 la_data_in[53]
port 97 nsew signal input
rlabel metal2 s 62384 0 62440 400 6 la_data_in[54]
port 98 nsew signal input
rlabel metal2 s 63392 0 63448 400 6 la_data_in[55]
port 99 nsew signal input
rlabel metal2 s 64400 0 64456 400 6 la_data_in[56]
port 100 nsew signal input
rlabel metal2 s 65408 0 65464 400 6 la_data_in[57]
port 101 nsew signal input
rlabel metal2 s 66416 0 66472 400 6 la_data_in[58]
port 102 nsew signal input
rlabel metal2 s 67424 0 67480 400 6 la_data_in[59]
port 103 nsew signal input
rlabel metal2 s 12992 0 13048 400 6 la_data_in[5]
port 104 nsew signal input
rlabel metal2 s 68432 0 68488 400 6 la_data_in[60]
port 105 nsew signal input
rlabel metal2 s 69440 0 69496 400 6 la_data_in[61]
port 106 nsew signal input
rlabel metal2 s 70448 0 70504 400 6 la_data_in[62]
port 107 nsew signal input
rlabel metal2 s 71456 0 71512 400 6 la_data_in[63]
port 108 nsew signal input
rlabel metal2 s 14000 0 14056 400 6 la_data_in[6]
port 109 nsew signal input
rlabel metal2 s 15008 0 15064 400 6 la_data_in[7]
port 110 nsew signal input
rlabel metal2 s 16016 0 16072 400 6 la_data_in[8]
port 111 nsew signal input
rlabel metal2 s 17024 0 17080 400 6 la_data_in[9]
port 112 nsew signal input
rlabel metal2 s 8288 0 8344 400 6 la_data_out[0]
port 113 nsew signal output
rlabel metal2 s 18368 0 18424 400 6 la_data_out[10]
port 114 nsew signal output
rlabel metal2 s 19376 0 19432 400 6 la_data_out[11]
port 115 nsew signal output
rlabel metal2 s 20384 0 20440 400 6 la_data_out[12]
port 116 nsew signal output
rlabel metal2 s 21392 0 21448 400 6 la_data_out[13]
port 117 nsew signal output
rlabel metal2 s 22400 0 22456 400 6 la_data_out[14]
port 118 nsew signal output
rlabel metal2 s 23408 0 23464 400 6 la_data_out[15]
port 119 nsew signal output
rlabel metal2 s 24416 0 24472 400 6 la_data_out[16]
port 120 nsew signal output
rlabel metal2 s 25424 0 25480 400 6 la_data_out[17]
port 121 nsew signal output
rlabel metal2 s 26432 0 26488 400 6 la_data_out[18]
port 122 nsew signal output
rlabel metal2 s 27440 0 27496 400 6 la_data_out[19]
port 123 nsew signal output
rlabel metal2 s 9296 0 9352 400 6 la_data_out[1]
port 124 nsew signal output
rlabel metal2 s 28448 0 28504 400 6 la_data_out[20]
port 125 nsew signal output
rlabel metal2 s 29456 0 29512 400 6 la_data_out[21]
port 126 nsew signal output
rlabel metal2 s 30464 0 30520 400 6 la_data_out[22]
port 127 nsew signal output
rlabel metal2 s 31472 0 31528 400 6 la_data_out[23]
port 128 nsew signal output
rlabel metal2 s 32480 0 32536 400 6 la_data_out[24]
port 129 nsew signal output
rlabel metal2 s 33488 0 33544 400 6 la_data_out[25]
port 130 nsew signal output
rlabel metal2 s 34496 0 34552 400 6 la_data_out[26]
port 131 nsew signal output
rlabel metal2 s 35504 0 35560 400 6 la_data_out[27]
port 132 nsew signal output
rlabel metal2 s 36512 0 36568 400 6 la_data_out[28]
port 133 nsew signal output
rlabel metal2 s 37520 0 37576 400 6 la_data_out[29]
port 134 nsew signal output
rlabel metal2 s 10304 0 10360 400 6 la_data_out[2]
port 135 nsew signal output
rlabel metal2 s 38528 0 38584 400 6 la_data_out[30]
port 136 nsew signal output
rlabel metal2 s 39536 0 39592 400 6 la_data_out[31]
port 137 nsew signal output
rlabel metal2 s 40544 0 40600 400 6 la_data_out[32]
port 138 nsew signal output
rlabel metal2 s 41552 0 41608 400 6 la_data_out[33]
port 139 nsew signal output
rlabel metal2 s 42560 0 42616 400 6 la_data_out[34]
port 140 nsew signal output
rlabel metal2 s 43568 0 43624 400 6 la_data_out[35]
port 141 nsew signal output
rlabel metal2 s 44576 0 44632 400 6 la_data_out[36]
port 142 nsew signal output
rlabel metal2 s 45584 0 45640 400 6 la_data_out[37]
port 143 nsew signal output
rlabel metal2 s 46592 0 46648 400 6 la_data_out[38]
port 144 nsew signal output
rlabel metal2 s 47600 0 47656 400 6 la_data_out[39]
port 145 nsew signal output
rlabel metal2 s 11312 0 11368 400 6 la_data_out[3]
port 146 nsew signal output
rlabel metal2 s 48608 0 48664 400 6 la_data_out[40]
port 147 nsew signal output
rlabel metal2 s 49616 0 49672 400 6 la_data_out[41]
port 148 nsew signal output
rlabel metal2 s 50624 0 50680 400 6 la_data_out[42]
port 149 nsew signal output
rlabel metal2 s 51632 0 51688 400 6 la_data_out[43]
port 150 nsew signal output
rlabel metal2 s 52640 0 52696 400 6 la_data_out[44]
port 151 nsew signal output
rlabel metal2 s 53648 0 53704 400 6 la_data_out[45]
port 152 nsew signal output
rlabel metal2 s 54656 0 54712 400 6 la_data_out[46]
port 153 nsew signal output
rlabel metal2 s 55664 0 55720 400 6 la_data_out[47]
port 154 nsew signal output
rlabel metal2 s 56672 0 56728 400 6 la_data_out[48]
port 155 nsew signal output
rlabel metal2 s 57680 0 57736 400 6 la_data_out[49]
port 156 nsew signal output
rlabel metal2 s 12320 0 12376 400 6 la_data_out[4]
port 157 nsew signal output
rlabel metal2 s 58688 0 58744 400 6 la_data_out[50]
port 158 nsew signal output
rlabel metal2 s 59696 0 59752 400 6 la_data_out[51]
port 159 nsew signal output
rlabel metal2 s 60704 0 60760 400 6 la_data_out[52]
port 160 nsew signal output
rlabel metal2 s 61712 0 61768 400 6 la_data_out[53]
port 161 nsew signal output
rlabel metal2 s 62720 0 62776 400 6 la_data_out[54]
port 162 nsew signal output
rlabel metal2 s 63728 0 63784 400 6 la_data_out[55]
port 163 nsew signal output
rlabel metal2 s 64736 0 64792 400 6 la_data_out[56]
port 164 nsew signal output
rlabel metal2 s 65744 0 65800 400 6 la_data_out[57]
port 165 nsew signal output
rlabel metal2 s 66752 0 66808 400 6 la_data_out[58]
port 166 nsew signal output
rlabel metal2 s 67760 0 67816 400 6 la_data_out[59]
port 167 nsew signal output
rlabel metal2 s 13328 0 13384 400 6 la_data_out[5]
port 168 nsew signal output
rlabel metal2 s 68768 0 68824 400 6 la_data_out[60]
port 169 nsew signal output
rlabel metal2 s 69776 0 69832 400 6 la_data_out[61]
port 170 nsew signal output
rlabel metal2 s 70784 0 70840 400 6 la_data_out[62]
port 171 nsew signal output
rlabel metal2 s 71792 0 71848 400 6 la_data_out[63]
port 172 nsew signal output
rlabel metal2 s 14336 0 14392 400 6 la_data_out[6]
port 173 nsew signal output
rlabel metal2 s 15344 0 15400 400 6 la_data_out[7]
port 174 nsew signal output
rlabel metal2 s 16352 0 16408 400 6 la_data_out[8]
port 175 nsew signal output
rlabel metal2 s 17360 0 17416 400 6 la_data_out[9]
port 176 nsew signal output
rlabel metal2 s 8624 0 8680 400 6 la_oenb[0]
port 177 nsew signal input
rlabel metal2 s 18704 0 18760 400 6 la_oenb[10]
port 178 nsew signal input
rlabel metal2 s 19712 0 19768 400 6 la_oenb[11]
port 179 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 la_oenb[12]
port 180 nsew signal input
rlabel metal2 s 21728 0 21784 400 6 la_oenb[13]
port 181 nsew signal input
rlabel metal2 s 22736 0 22792 400 6 la_oenb[14]
port 182 nsew signal input
rlabel metal2 s 23744 0 23800 400 6 la_oenb[15]
port 183 nsew signal input
rlabel metal2 s 24752 0 24808 400 6 la_oenb[16]
port 184 nsew signal input
rlabel metal2 s 25760 0 25816 400 6 la_oenb[17]
port 185 nsew signal input
rlabel metal2 s 26768 0 26824 400 6 la_oenb[18]
port 186 nsew signal input
rlabel metal2 s 27776 0 27832 400 6 la_oenb[19]
port 187 nsew signal input
rlabel metal2 s 9632 0 9688 400 6 la_oenb[1]
port 188 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 la_oenb[20]
port 189 nsew signal input
rlabel metal2 s 29792 0 29848 400 6 la_oenb[21]
port 190 nsew signal input
rlabel metal2 s 30800 0 30856 400 6 la_oenb[22]
port 191 nsew signal input
rlabel metal2 s 31808 0 31864 400 6 la_oenb[23]
port 192 nsew signal input
rlabel metal2 s 32816 0 32872 400 6 la_oenb[24]
port 193 nsew signal input
rlabel metal2 s 33824 0 33880 400 6 la_oenb[25]
port 194 nsew signal input
rlabel metal2 s 34832 0 34888 400 6 la_oenb[26]
port 195 nsew signal input
rlabel metal2 s 35840 0 35896 400 6 la_oenb[27]
port 196 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 la_oenb[28]
port 197 nsew signal input
rlabel metal2 s 37856 0 37912 400 6 la_oenb[29]
port 198 nsew signal input
rlabel metal2 s 10640 0 10696 400 6 la_oenb[2]
port 199 nsew signal input
rlabel metal2 s 38864 0 38920 400 6 la_oenb[30]
port 200 nsew signal input
rlabel metal2 s 39872 0 39928 400 6 la_oenb[31]
port 201 nsew signal input
rlabel metal2 s 40880 0 40936 400 6 la_oenb[32]
port 202 nsew signal input
rlabel metal2 s 41888 0 41944 400 6 la_oenb[33]
port 203 nsew signal input
rlabel metal2 s 42896 0 42952 400 6 la_oenb[34]
port 204 nsew signal input
rlabel metal2 s 43904 0 43960 400 6 la_oenb[35]
port 205 nsew signal input
rlabel metal2 s 44912 0 44968 400 6 la_oenb[36]
port 206 nsew signal input
rlabel metal2 s 45920 0 45976 400 6 la_oenb[37]
port 207 nsew signal input
rlabel metal2 s 46928 0 46984 400 6 la_oenb[38]
port 208 nsew signal input
rlabel metal2 s 47936 0 47992 400 6 la_oenb[39]
port 209 nsew signal input
rlabel metal2 s 11648 0 11704 400 6 la_oenb[3]
port 210 nsew signal input
rlabel metal2 s 48944 0 49000 400 6 la_oenb[40]
port 211 nsew signal input
rlabel metal2 s 49952 0 50008 400 6 la_oenb[41]
port 212 nsew signal input
rlabel metal2 s 50960 0 51016 400 6 la_oenb[42]
port 213 nsew signal input
rlabel metal2 s 51968 0 52024 400 6 la_oenb[43]
port 214 nsew signal input
rlabel metal2 s 52976 0 53032 400 6 la_oenb[44]
port 215 nsew signal input
rlabel metal2 s 53984 0 54040 400 6 la_oenb[45]
port 216 nsew signal input
rlabel metal2 s 54992 0 55048 400 6 la_oenb[46]
port 217 nsew signal input
rlabel metal2 s 56000 0 56056 400 6 la_oenb[47]
port 218 nsew signal input
rlabel metal2 s 57008 0 57064 400 6 la_oenb[48]
port 219 nsew signal input
rlabel metal2 s 58016 0 58072 400 6 la_oenb[49]
port 220 nsew signal input
rlabel metal2 s 12656 0 12712 400 6 la_oenb[4]
port 221 nsew signal input
rlabel metal2 s 59024 0 59080 400 6 la_oenb[50]
port 222 nsew signal input
rlabel metal2 s 60032 0 60088 400 6 la_oenb[51]
port 223 nsew signal input
rlabel metal2 s 61040 0 61096 400 6 la_oenb[52]
port 224 nsew signal input
rlabel metal2 s 62048 0 62104 400 6 la_oenb[53]
port 225 nsew signal input
rlabel metal2 s 63056 0 63112 400 6 la_oenb[54]
port 226 nsew signal input
rlabel metal2 s 64064 0 64120 400 6 la_oenb[55]
port 227 nsew signal input
rlabel metal2 s 65072 0 65128 400 6 la_oenb[56]
port 228 nsew signal input
rlabel metal2 s 66080 0 66136 400 6 la_oenb[57]
port 229 nsew signal input
rlabel metal2 s 67088 0 67144 400 6 la_oenb[58]
port 230 nsew signal input
rlabel metal2 s 68096 0 68152 400 6 la_oenb[59]
port 231 nsew signal input
rlabel metal2 s 13664 0 13720 400 6 la_oenb[5]
port 232 nsew signal input
rlabel metal2 s 69104 0 69160 400 6 la_oenb[60]
port 233 nsew signal input
rlabel metal2 s 70112 0 70168 400 6 la_oenb[61]
port 234 nsew signal input
rlabel metal2 s 71120 0 71176 400 6 la_oenb[62]
port 235 nsew signal input
rlabel metal2 s 72128 0 72184 400 6 la_oenb[63]
port 236 nsew signal input
rlabel metal2 s 14672 0 14728 400 6 la_oenb[6]
port 237 nsew signal input
rlabel metal2 s 15680 0 15736 400 6 la_oenb[7]
port 238 nsew signal input
rlabel metal2 s 16688 0 16744 400 6 la_oenb[8]
port 239 nsew signal input
rlabel metal2 s 17696 0 17752 400 6 la_oenb[9]
port 240 nsew signal input
rlabel metal4 s 2224 1538 2384 78430 6 vdd
port 241 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 78430 6 vdd
port 241 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 78430 6 vdd
port 241 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 78430 6 vdd
port 241 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 78430 6 vdd
port 241 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 78430 6 vdd
port 241 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 78430 6 vss
port 242 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 78430 6 vss
port 242 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 78430 6 vss
port 242 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 78430 6 vss
port 242 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 78430 6 vss
port 242 nsew ground bidirectional
rlabel metal2 s 7616 0 7672 400 6 wb_clk_i
port 243 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 80000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12848914
string GDS_FILE /home/kris/repos/diy-ic/lincoln-gfmpw-1d/openlane/user_proj_example/runs/23_12_08_02_22/results/signoff/user_proj_example.magic.gds
string GDS_START 383064
<< end >>

