magic
tech gf180mcuD
magscale 1 5
timestamp 1701888964
<< obsm1 >>
rect 672 1538 77056 77769
<< metal2 >>
rect 47712 79134 47768 79534
rect 48048 79134 48104 79534
rect 48384 79134 48440 79534
rect 48720 79134 48776 79534
rect 49056 79134 49112 79534
rect 49392 79134 49448 79534
rect 49728 79134 49784 79534
rect 50064 79134 50120 79534
rect 50400 79134 50456 79534
rect 50736 79134 50792 79534
rect 51072 79134 51128 79534
rect 52080 79134 52136 79534
rect 28560 0 28616 400
rect 28896 0 28952 400
rect 29232 0 29288 400
rect 29904 0 29960 400
rect 30240 0 30296 400
rect 30576 0 30632 400
rect 30912 0 30968 400
rect 31248 0 31304 400
rect 32256 0 32312 400
rect 32928 0 32984 400
rect 33264 0 33320 400
rect 33936 0 33992 400
rect 36288 0 36344 400
rect 36624 0 36680 400
rect 36960 0 37016 400
rect 49392 0 49448 400
rect 49728 0 49784 400
rect 50064 0 50120 400
rect 50400 0 50456 400
rect 67200 0 67256 400
rect 67536 0 67592 400
rect 67872 0 67928 400
rect 68208 0 68264 400
rect 68544 0 68600 400
rect 68880 0 68936 400
<< obsm2 >>
rect 14 79104 47682 79134
rect 47798 79104 48018 79134
rect 48134 79104 48354 79134
rect 48470 79104 48690 79134
rect 48806 79104 49026 79134
rect 49142 79104 49362 79134
rect 49478 79104 49698 79134
rect 49814 79104 50034 79134
rect 50150 79104 50370 79134
rect 50486 79104 50706 79134
rect 50822 79104 51042 79134
rect 51158 79104 52050 79134
rect 52166 79104 76874 79134
rect 14 430 76874 79104
rect 14 350 28530 430
rect 28646 350 28866 430
rect 28982 350 29202 430
rect 29318 350 29874 430
rect 29990 350 30210 430
rect 30326 350 30546 430
rect 30662 350 30882 430
rect 30998 350 31218 430
rect 31334 350 32226 430
rect 32342 350 32898 430
rect 33014 350 33234 430
rect 33350 350 33906 430
rect 34022 350 36258 430
rect 36374 350 36594 430
rect 36710 350 36930 430
rect 37046 350 49362 430
rect 49478 350 49698 430
rect 49814 350 50034 430
rect 50150 350 50370 430
rect 50486 350 67170 430
rect 67286 350 67506 430
rect 67622 350 67842 430
rect 67958 350 68178 430
rect 68294 350 68514 430
rect 68630 350 68850 430
rect 68966 350 76874 430
<< metal3 >>
rect 0 76608 400 76664
rect 0 57456 400 57512
rect 0 57120 400 57176
rect 0 56784 400 56840
rect 0 55440 400 55496
rect 0 54432 400 54488
rect 0 53424 400 53480
rect 0 52080 400 52136
rect 0 50400 400 50456
rect 0 49392 400 49448
rect 0 49056 400 49112
rect 0 48720 400 48776
rect 0 48384 400 48440
rect 0 48048 400 48104
rect 0 47712 400 47768
rect 77342 47712 77742 47768
rect 0 47376 400 47432
rect 77342 47376 77742 47432
rect 0 47040 400 47096
rect 0 46704 400 46760
rect 0 46368 400 46424
rect 0 46032 400 46088
rect 77342 46032 77742 46088
rect 0 45696 400 45752
rect 77342 45696 77742 45752
rect 77342 45024 77742 45080
rect 77342 44352 77742 44408
rect 77342 44016 77742 44072
rect 77342 43344 77742 43400
rect 77342 42672 77742 42728
rect 77342 32256 77742 32312
rect 0 26544 400 26600
rect 0 26208 400 26264
rect 77342 23184 77742 23240
rect 0 12096 400 12152
<< obsm3 >>
rect 9 76694 77342 77630
rect 430 76578 77342 76694
rect 9 57542 77342 76578
rect 430 57426 77342 57542
rect 9 57206 77342 57426
rect 430 57090 77342 57206
rect 9 56870 77342 57090
rect 430 56754 77342 56870
rect 9 55526 77342 56754
rect 430 55410 77342 55526
rect 9 54518 77342 55410
rect 430 54402 77342 54518
rect 9 53510 77342 54402
rect 430 53394 77342 53510
rect 9 52166 77342 53394
rect 430 52050 77342 52166
rect 9 50486 77342 52050
rect 430 50370 77342 50486
rect 9 49478 77342 50370
rect 430 49362 77342 49478
rect 9 49142 77342 49362
rect 430 49026 77342 49142
rect 9 48806 77342 49026
rect 430 48690 77342 48806
rect 9 48470 77342 48690
rect 430 48354 77342 48470
rect 9 48134 77342 48354
rect 430 48018 77342 48134
rect 9 47798 77342 48018
rect 430 47682 77312 47798
rect 9 47462 77342 47682
rect 430 47346 77312 47462
rect 9 47126 77342 47346
rect 430 47010 77342 47126
rect 9 46790 77342 47010
rect 430 46674 77342 46790
rect 9 46454 77342 46674
rect 430 46338 77342 46454
rect 9 46118 77342 46338
rect 430 46002 77312 46118
rect 9 45782 77342 46002
rect 430 45666 77312 45782
rect 9 45110 77342 45666
rect 9 44994 77312 45110
rect 9 44438 77342 44994
rect 9 44322 77312 44438
rect 9 44102 77342 44322
rect 9 43986 77312 44102
rect 9 43430 77342 43986
rect 9 43314 77312 43430
rect 9 42758 77342 43314
rect 9 42642 77312 42758
rect 9 32342 77342 42642
rect 9 32226 77312 32342
rect 9 26630 77342 32226
rect 430 26514 77342 26630
rect 9 26294 77342 26514
rect 430 26178 77342 26294
rect 9 23270 77342 26178
rect 9 23154 77312 23270
rect 9 12182 77342 23154
rect 430 12066 77342 12182
rect 9 630 77342 12066
<< metal4 >>
rect 2224 1538 2384 77646
rect 9904 1538 10064 77646
rect 17584 1538 17744 77646
rect 25264 1538 25424 77646
rect 32944 1538 33104 77646
rect 40624 1538 40784 77646
rect 48304 1538 48464 77646
rect 55984 1538 56144 77646
rect 63664 1538 63824 77646
rect 71344 1538 71504 77646
<< obsm4 >>
rect 5670 1689 9874 77383
rect 10094 1689 17554 77383
rect 17774 1689 25234 77383
rect 25454 1689 32914 77383
rect 33134 1689 40594 77383
rect 40814 1689 48274 77383
rect 48494 1689 55954 77383
rect 56174 1689 63634 77383
rect 63854 1689 71314 77383
rect 71534 1689 72226 77383
<< labels >>
rlabel metal3 s 77342 44016 77742 44072 6 address_i[0]
port 1 nsew signal input
rlabel metal3 s 77342 23184 77742 23240 6 address_i[1]
port 2 nsew signal input
rlabel metal3 s 77342 32256 77742 32312 6 address_i[2]
port 3 nsew signal input
rlabel metal2 s 36288 0 36344 400 6 address_i[3]
port 4 nsew signal input
rlabel metal2 s 36624 0 36680 400 6 address_i[4]
port 5 nsew signal input
rlabel metal2 s 36960 0 37016 400 6 address_i[5]
port 6 nsew signal input
rlabel metal3 s 0 76608 400 76664 6 clk_i
port 7 nsew signal input
rlabel metal2 s 33936 0 33992 400 6 data_i[0]
port 8 nsew signal input
rlabel metal3 s 77342 42672 77742 42728 6 data_i[10]
port 9 nsew signal input
rlabel metal3 s 77342 43344 77742 43400 6 data_i[11]
port 10 nsew signal input
rlabel metal3 s 77342 44352 77742 44408 6 data_i[12]
port 11 nsew signal input
rlabel metal3 s 77342 45024 77742 45080 6 data_i[13]
port 12 nsew signal input
rlabel metal2 s 48720 79134 48776 79534 6 data_i[14]
port 13 nsew signal input
rlabel metal2 s 47712 79134 47768 79534 6 data_i[15]
port 14 nsew signal input
rlabel metal2 s 48048 79134 48104 79534 6 data_i[16]
port 15 nsew signal input
rlabel metal2 s 48384 79134 48440 79534 6 data_i[17]
port 16 nsew signal input
rlabel metal2 s 49056 79134 49112 79534 6 data_i[18]
port 17 nsew signal input
rlabel metal2 s 49392 79134 49448 79534 6 data_i[19]
port 18 nsew signal input
rlabel metal2 s 32928 0 32984 400 6 data_i[1]
port 19 nsew signal input
rlabel metal3 s 0 45696 400 45752 6 data_i[20]
port 20 nsew signal input
rlabel metal3 s 0 46032 400 46088 6 data_i[21]
port 21 nsew signal input
rlabel metal3 s 0 48384 400 48440 6 data_i[22]
port 22 nsew signal input
rlabel metal3 s 0 46368 400 46424 6 data_i[23]
port 23 nsew signal input
rlabel metal3 s 0 47040 400 47096 6 data_i[24]
port 24 nsew signal input
rlabel metal3 s 0 47376 400 47432 6 data_i[25]
port 25 nsew signal input
rlabel metal3 s 0 49056 400 49112 6 data_i[26]
port 26 nsew signal input
rlabel metal3 s 0 48048 400 48104 6 data_i[27]
port 27 nsew signal input
rlabel metal3 s 0 46704 400 46760 6 data_i[28]
port 28 nsew signal input
rlabel metal3 s 0 48720 400 48776 6 data_i[29]
port 29 nsew signal input
rlabel metal2 s 31248 0 31304 400 6 data_i[2]
port 30 nsew signal input
rlabel metal2 s 28560 0 28616 400 6 data_i[30]
port 31 nsew signal input
rlabel metal2 s 28896 0 28952 400 6 data_i[31]
port 32 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 data_i[3]
port 33 nsew signal input
rlabel metal2 s 32256 0 32312 400 6 data_i[4]
port 34 nsew signal input
rlabel metal2 s 30576 0 30632 400 6 data_i[5]
port 35 nsew signal input
rlabel metal2 s 30912 0 30968 400 6 data_i[6]
port 36 nsew signal input
rlabel metal2 s 29904 0 29960 400 6 data_i[7]
port 37 nsew signal input
rlabel metal2 s 29232 0 29288 400 6 data_i[8]
port 38 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 data_i[9]
port 39 nsew signal input
rlabel metal2 s 49728 0 49784 400 6 data_o[0]
port 40 nsew signal output
rlabel metal3 s 77342 46032 77742 46088 6 data_o[10]
port 41 nsew signal output
rlabel metal2 s 50736 79134 50792 79534 6 data_o[11]
port 42 nsew signal output
rlabel metal3 s 77342 45696 77742 45752 6 data_o[12]
port 43 nsew signal output
rlabel metal2 s 50400 79134 50456 79534 6 data_o[13]
port 44 nsew signal output
rlabel metal3 s 77342 47712 77742 47768 6 data_o[14]
port 45 nsew signal output
rlabel metal3 s 77342 47376 77742 47432 6 data_o[15]
port 46 nsew signal output
rlabel metal2 s 52080 79134 52136 79534 6 data_o[16]
port 47 nsew signal output
rlabel metal2 s 50064 79134 50120 79534 6 data_o[17]
port 48 nsew signal output
rlabel metal2 s 51072 79134 51128 79534 6 data_o[18]
port 49 nsew signal output
rlabel metal2 s 49728 79134 49784 79534 6 data_o[19]
port 50 nsew signal output
rlabel metal2 s 49392 0 49448 400 6 data_o[1]
port 51 nsew signal output
rlabel metal3 s 0 57120 400 57176 6 data_o[20]
port 52 nsew signal output
rlabel metal3 s 0 57456 400 57512 6 data_o[21]
port 53 nsew signal output
rlabel metal3 s 0 55440 400 55496 6 data_o[22]
port 54 nsew signal output
rlabel metal3 s 0 56784 400 56840 6 data_o[23]
port 55 nsew signal output
rlabel metal3 s 0 53424 400 53480 6 data_o[24]
port 56 nsew signal output
rlabel metal3 s 0 54432 400 54488 6 data_o[25]
port 57 nsew signal output
rlabel metal3 s 0 52080 400 52136 6 data_o[26]
port 58 nsew signal output
rlabel metal3 s 0 50400 400 50456 6 data_o[27]
port 59 nsew signal output
rlabel metal3 s 0 49392 400 49448 6 data_o[28]
port 60 nsew signal output
rlabel metal3 s 0 47712 400 47768 6 data_o[29]
port 61 nsew signal output
rlabel metal2 s 50064 0 50120 400 6 data_o[2]
port 62 nsew signal output
rlabel metal3 s 0 26544 400 26600 6 data_o[30]
port 63 nsew signal output
rlabel metal3 s 0 26208 400 26264 6 data_o[31]
port 64 nsew signal output
rlabel metal2 s 50400 0 50456 400 6 data_o[3]
port 65 nsew signal output
rlabel metal2 s 68880 0 68936 400 6 data_o[4]
port 66 nsew signal output
rlabel metal2 s 67536 0 67592 400 6 data_o[5]
port 67 nsew signal output
rlabel metal2 s 68208 0 68264 400 6 data_o[6]
port 68 nsew signal output
rlabel metal2 s 67872 0 67928 400 6 data_o[7]
port 69 nsew signal output
rlabel metal2 s 67200 0 67256 400 6 data_o[8]
port 70 nsew signal output
rlabel metal2 s 68544 0 68600 400 6 data_o[9]
port 71 nsew signal output
rlabel metal4 s 2224 1538 2384 77646 6 vdd
port 72 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 77646 6 vdd
port 72 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 77646 6 vdd
port 72 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 77646 6 vdd
port 72 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 77646 6 vdd
port 72 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 77646 6 vss
port 73 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 77646 6 vss
port 73 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 77646 6 vss
port 73 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 77646 6 vss
port 73 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 77646 6 vss
port 73 nsew ground bidirectional
rlabel metal3 s 0 12096 400 12152 6 we_i
port 74 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 77742 79534
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 18575976
string GDS_FILE /home/kris/repos/diy-ic/lincoln-gfmpw/openlane/ram_6x64/runs/23_12_06_18_46/results/signoff/ram_6x64.magic.gds
string GDS_START 248100
<< end >>

