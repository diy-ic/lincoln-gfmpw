VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO titan
  CLASS BLOCK ;
  FOREIGN titan ;
  ORIGIN 0.000 0.000 ;
  SIZE 586.805 BY 604.725 ;
  PIN spi_clock_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 0.000 276.080 4.000 ;
    END
  END spi_clock_i
  PIN spi_cs_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 0.000 279.440 4.000 ;
    END
  END spi_cs_i
  PIN spi_pico_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 0.000 353.360 4.000 ;
    END
  END spi_pico_i
  PIN spi_poci_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 0.000 306.320 4.000 ;
    END
  END spi_poci_o
  PIN sys_clock_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 561.120 4.000 561.680 ;
    END
  END sys_clock_i
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 588.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 588.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 588.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 588.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 588.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 588.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 588.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 588.300 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 579.600 588.300 ;
      LAYER Metal2 ;
        RECT 9.660 4.300 577.780 588.190 ;
        RECT 9.660 4.000 275.220 4.300 ;
        RECT 276.380 4.000 278.580 4.300 ;
        RECT 279.740 4.000 305.460 4.300 ;
        RECT 306.620 4.000 352.500 4.300 ;
        RECT 353.660 4.000 577.780 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 561.980 577.830 588.140 ;
        RECT 4.300 560.820 577.830 561.980 ;
        RECT 4.000 15.540 577.830 560.820 ;
      LAYER Metal4 ;
        RECT 15.260 33.690 21.940 572.790 ;
        RECT 24.140 33.690 98.740 572.790 ;
        RECT 100.940 33.690 175.540 572.790 ;
        RECT 177.740 33.690 252.340 572.790 ;
        RECT 254.540 33.690 329.140 572.790 ;
        RECT 331.340 33.690 405.940 572.790 ;
        RECT 408.140 33.690 482.740 572.790 ;
        RECT 484.940 33.690 544.740 572.790 ;
  END
END titan
END LIBRARY

