VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO titan
  CLASS BLOCK ;
  FOREIGN titan ;
  ORIGIN 0.000 0.000 ;
  SIZE 526.275 BY 544.195 ;
  PIN spi_clock_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 0.000 259.280 4.000 ;
    END
  END spi_clock_i
  PIN spi_cs_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 0.000 262.640 4.000 ;
    END
  END spi_cs_i
  PIN spi_pico_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 0.000 339.920 4.000 ;
    END
  END spi_pico_i
  PIN spi_poci_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 0.000 289.520 4.000 ;
    END
  END spi_poci_o
  PIN sys_clock_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 517.440 4.000 518.000 ;
    END
  END sys_clock_i
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 525.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 525.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 525.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 525.580 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 525.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 525.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 525.580 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 519.120 526.250 ;
      LAYER Metal2 ;
        RECT 6.300 4.300 516.740 526.310 ;
        RECT 6.300 4.000 258.420 4.300 ;
        RECT 259.580 4.000 261.780 4.300 ;
        RECT 262.940 4.000 288.660 4.300 ;
        RECT 289.820 4.000 339.060 4.300 ;
        RECT 340.220 4.000 516.740 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 518.300 516.790 525.420 ;
        RECT 4.300 517.140 516.790 518.300 ;
        RECT 4.000 15.540 516.790 517.140 ;
      LAYER Metal4 ;
        RECT 16.940 21.930 21.940 477.590 ;
        RECT 24.140 21.930 98.740 477.590 ;
        RECT 100.940 21.930 175.540 477.590 ;
        RECT 177.740 21.930 252.340 477.590 ;
        RECT 254.540 21.930 329.140 477.590 ;
        RECT 331.340 21.930 405.940 477.590 ;
        RECT 408.140 21.930 482.740 477.590 ;
        RECT 484.940 21.930 487.060 477.590 ;
  END
END titan
END LIBRARY

