VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ram
  CLASS BLOCK ;
  FOREIGN ram ;
  ORIGIN 0.000 0.000 ;
  SIZE 556.985 BY 574.905 ;
  PIN address_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 312.480 4.000 313.040 ;
    END
  END address_i[0]
  PIN address_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 292.320 4.000 292.880 ;
    END
  END address_i[1]
  PIN address_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.600 4.000 286.160 ;
    END
  END address_i[2]
  PIN address_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 285.600 556.985 286.160 ;
    END
  END address_i[3]
  PIN address_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 0.000 306.320 4.000 ;
    END
  END address_i[4]
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 547.680 4.000 548.240 ;
    END
  END clk_i
  PIN data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 258.720 556.985 259.280 ;
    END
  END data_i[0]
  PIN data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 570.905 319.760 574.905 ;
    END
  END data_i[10]
  PIN data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 570.905 323.120 574.905 ;
    END
  END data_i[11]
  PIN data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 570.905 306.320 574.905 ;
    END
  END data_i[12]
  PIN data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 570.905 279.440 574.905 ;
    END
  END data_i[13]
  PIN data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 570.905 262.640 574.905 ;
    END
  END data_i[14]
  PIN data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 570.905 235.760 574.905 ;
    END
  END data_i[15]
  PIN data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 570.905 239.120 574.905 ;
    END
  END data_i[16]
  PIN data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 570.905 232.400 574.905 ;
    END
  END data_i[17]
  PIN data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 570.905 252.560 574.905 ;
    END
  END data_i[18]
  PIN data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 570.905 242.480 574.905 ;
    END
  END data_i[19]
  PIN data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 262.080 556.985 262.640 ;
    END
  END data_i[1]
  PIN data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 0.000 239.120 4.000 ;
    END
  END data_i[20]
  PIN data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 4.000 ;
    END
  END data_i[21]
  PIN data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END data_i[22]
  PIN data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 4.000 145.040 ;
    END
  END data_i[23]
  PIN data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END data_i[24]
  PIN data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END data_i[25]
  PIN data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END data_i[26]
  PIN data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 4.000 158.480 ;
    END
  END data_i[27]
  PIN data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 0.000 235.760 4.000 ;
    END
  END data_i[28]
  PIN data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 0.000 269.360 4.000 ;
    END
  END data_i[29]
  PIN data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 265.440 556.985 266.000 ;
    END
  END data_i[2]
  PIN data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 0.000 276.080 4.000 ;
    END
  END data_i[30]
  PIN data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 0.000 316.400 4.000 ;
    END
  END data_i[31]
  PIN data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 288.960 556.985 289.520 ;
    END
  END data_i[3]
  PIN data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 312.480 556.985 313.040 ;
    END
  END data_i[4]
  PIN data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 356.160 556.985 356.720 ;
    END
  END data_i[5]
  PIN data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 393.120 556.985 393.680 ;
    END
  END data_i[6]
  PIN data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 409.920 556.985 410.480 ;
    END
  END data_i[7]
  PIN data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 396.480 556.985 397.040 ;
    END
  END data_i[8]
  PIN data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 570.905 343.280 574.905 ;
    END
  END data_i[9]
  PIN data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 211.680 556.985 212.240 ;
    END
  END data_o[0]
  PIN data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 570.905 192.080 574.905 ;
    END
  END data_o[10]
  PIN data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 570.905 188.720 574.905 ;
    END
  END data_o[11]
  PIN data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 570.905 185.360 574.905 ;
    END
  END data_o[12]
  PIN data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 570.905 171.920 574.905 ;
    END
  END data_o[13]
  PIN data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 570.905 168.560 574.905 ;
    END
  END data_o[14]
  PIN data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 570.905 165.200 574.905 ;
    END
  END data_o[15]
  PIN data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 570.905 195.440 574.905 ;
    END
  END data_o[16]
  PIN data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 396.480 4.000 397.040 ;
    END
  END data_o[17]
  PIN data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 352.800 4.000 353.360 ;
    END
  END data_o[18]
  PIN data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.720 4.000 343.280 ;
    END
  END data_o[19]
  PIN data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 215.040 556.985 215.600 ;
    END
  END data_o[1]
  PIN data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 0.000 175.280 4.000 ;
    END
  END data_o[20]
  PIN data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 181.440 4.000 182.000 ;
    END
  END data_o[21]
  PIN data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END data_o[22]
  PIN data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.720 4.000 175.280 ;
    END
  END data_o[23]
  PIN data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 171.360 4.000 171.920 ;
    END
  END data_o[24]
  PIN data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.160 4.000 188.720 ;
    END
  END data_o[25]
  PIN data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 4.000 195.440 ;
    END
  END data_o[26]
  PIN data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END data_o[27]
  PIN data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 4.000 185.360 ;
    END
  END data_o[28]
  PIN data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.520 4.000 192.080 ;
    END
  END data_o[29]
  PIN data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 208.320 556.985 208.880 ;
    END
  END data_o[2]
  PIN data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 0.000 323.120 4.000 ;
    END
  END data_o[30]
  PIN data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 0.000 350.000 4.000 ;
    END
  END data_o[31]
  PIN data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 241.920 556.985 242.480 ;
    END
  END data_o[3]
  PIN data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 315.840 556.985 316.400 ;
    END
  END data_o[4]
  PIN data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 322.560 556.985 323.120 ;
    END
  END data_o[5]
  PIN data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 336.000 556.985 336.560 ;
    END
  END data_o[6]
  PIN data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 332.640 556.985 333.200 ;
    END
  END data_o[7]
  PIN data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 346.080 556.985 346.640 ;
    END
  END data_o[8]
  PIN data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 552.985 352.800 556.985 353.360 ;
    END
  END data_o[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 556.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 556.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 556.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 556.940 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 556.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 556.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 556.940 ;
    END
  END vss
  PIN we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 299.040 4.000 299.600 ;
    END
  END we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 549.920 558.730 ;
      LAYER Metal2 ;
        RECT 8.540 570.605 164.340 570.905 ;
        RECT 165.500 570.605 167.700 570.905 ;
        RECT 168.860 570.605 171.060 570.905 ;
        RECT 172.220 570.605 184.500 570.905 ;
        RECT 185.660 570.605 187.860 570.905 ;
        RECT 189.020 570.605 191.220 570.905 ;
        RECT 192.380 570.605 194.580 570.905 ;
        RECT 195.740 570.605 231.540 570.905 ;
        RECT 232.700 570.605 234.900 570.905 ;
        RECT 236.060 570.605 238.260 570.905 ;
        RECT 239.420 570.605 241.620 570.905 ;
        RECT 242.780 570.605 251.700 570.905 ;
        RECT 252.860 570.605 261.780 570.905 ;
        RECT 262.940 570.605 278.580 570.905 ;
        RECT 279.740 570.605 305.460 570.905 ;
        RECT 306.620 570.605 318.900 570.905 ;
        RECT 320.060 570.605 322.260 570.905 ;
        RECT 323.420 570.605 342.420 570.905 ;
        RECT 343.580 570.605 553.700 570.905 ;
        RECT 8.540 4.300 553.700 570.605 ;
        RECT 8.540 3.500 110.580 4.300 ;
        RECT 111.740 3.500 160.980 4.300 ;
        RECT 162.140 3.500 167.700 4.300 ;
        RECT 168.860 3.500 174.420 4.300 ;
        RECT 175.580 3.500 177.780 4.300 ;
        RECT 178.940 3.500 234.900 4.300 ;
        RECT 236.060 3.500 238.260 4.300 ;
        RECT 239.420 3.500 268.500 4.300 ;
        RECT 269.660 3.500 275.220 4.300 ;
        RECT 276.380 3.500 305.460 4.300 ;
        RECT 306.620 3.500 315.540 4.300 ;
        RECT 316.700 3.500 322.260 4.300 ;
        RECT 323.420 3.500 349.140 4.300 ;
        RECT 350.300 3.500 553.700 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 548.540 553.700 562.660 ;
        RECT 4.300 547.380 553.700 548.540 ;
        RECT 4.000 410.780 553.700 547.380 ;
        RECT 4.000 409.620 552.685 410.780 ;
        RECT 4.000 397.340 553.700 409.620 ;
        RECT 4.300 396.180 552.685 397.340 ;
        RECT 4.000 393.980 553.700 396.180 ;
        RECT 4.000 392.820 552.685 393.980 ;
        RECT 4.000 357.020 553.700 392.820 ;
        RECT 4.000 355.860 552.685 357.020 ;
        RECT 4.000 353.660 553.700 355.860 ;
        RECT 4.300 352.500 552.685 353.660 ;
        RECT 4.000 346.940 553.700 352.500 ;
        RECT 4.000 345.780 552.685 346.940 ;
        RECT 4.000 343.580 553.700 345.780 ;
        RECT 4.300 342.420 553.700 343.580 ;
        RECT 4.000 336.860 553.700 342.420 ;
        RECT 4.000 335.700 552.685 336.860 ;
        RECT 4.000 333.500 553.700 335.700 ;
        RECT 4.000 332.340 552.685 333.500 ;
        RECT 4.000 323.420 553.700 332.340 ;
        RECT 4.000 322.260 552.685 323.420 ;
        RECT 4.000 316.700 553.700 322.260 ;
        RECT 4.000 315.540 552.685 316.700 ;
        RECT 4.000 313.340 553.700 315.540 ;
        RECT 4.300 312.180 552.685 313.340 ;
        RECT 4.000 299.900 553.700 312.180 ;
        RECT 4.300 298.740 553.700 299.900 ;
        RECT 4.000 293.180 553.700 298.740 ;
        RECT 4.300 292.020 553.700 293.180 ;
        RECT 4.000 289.820 553.700 292.020 ;
        RECT 4.000 288.660 552.685 289.820 ;
        RECT 4.000 286.460 553.700 288.660 ;
        RECT 4.300 285.300 552.685 286.460 ;
        RECT 4.000 266.300 553.700 285.300 ;
        RECT 4.000 265.140 552.685 266.300 ;
        RECT 4.000 262.940 553.700 265.140 ;
        RECT 4.000 261.780 552.685 262.940 ;
        RECT 4.000 259.580 553.700 261.780 ;
        RECT 4.000 258.420 552.685 259.580 ;
        RECT 4.000 242.780 553.700 258.420 ;
        RECT 4.000 241.620 552.685 242.780 ;
        RECT 4.000 215.900 553.700 241.620 ;
        RECT 4.000 214.740 552.685 215.900 ;
        RECT 4.000 212.540 553.700 214.740 ;
        RECT 4.000 211.380 552.685 212.540 ;
        RECT 4.000 209.180 553.700 211.380 ;
        RECT 4.000 208.020 552.685 209.180 ;
        RECT 4.000 195.740 553.700 208.020 ;
        RECT 4.300 194.580 553.700 195.740 ;
        RECT 4.000 192.380 553.700 194.580 ;
        RECT 4.300 191.220 553.700 192.380 ;
        RECT 4.000 189.020 553.700 191.220 ;
        RECT 4.300 187.860 553.700 189.020 ;
        RECT 4.000 185.660 553.700 187.860 ;
        RECT 4.300 184.500 553.700 185.660 ;
        RECT 4.000 182.300 553.700 184.500 ;
        RECT 4.300 181.140 553.700 182.300 ;
        RECT 4.000 175.580 553.700 181.140 ;
        RECT 4.300 174.420 553.700 175.580 ;
        RECT 4.000 172.220 553.700 174.420 ;
        RECT 4.300 171.060 553.700 172.220 ;
        RECT 4.000 168.860 553.700 171.060 ;
        RECT 4.300 167.700 553.700 168.860 ;
        RECT 4.000 158.780 553.700 167.700 ;
        RECT 4.300 157.620 553.700 158.780 ;
        RECT 4.000 145.340 553.700 157.620 ;
        RECT 4.300 144.180 553.700 145.340 ;
        RECT 4.000 128.540 553.700 144.180 ;
        RECT 4.300 127.380 553.700 128.540 ;
        RECT 4.000 115.100 553.700 127.380 ;
        RECT 4.300 113.940 553.700 115.100 ;
        RECT 4.000 15.540 553.700 113.940 ;
      LAYER Metal4 ;
        RECT 9.660 16.330 21.940 554.870 ;
        RECT 24.140 16.330 98.740 554.870 ;
        RECT 100.940 16.330 175.540 554.870 ;
        RECT 177.740 16.330 252.340 554.870 ;
        RECT 254.540 16.330 329.140 554.870 ;
        RECT 331.340 16.330 405.940 554.870 ;
        RECT 408.140 16.330 482.740 554.870 ;
        RECT 484.940 16.330 547.540 554.870 ;
  END
END ram
END LIBRARY

