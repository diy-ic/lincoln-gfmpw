magic
tech gf180mcuD
magscale 1 5
timestamp 1702036634
<< obsm1 >>
rect 672 1538 51912 52625
<< metal2 >>
rect 25872 0 25928 400
rect 26208 0 26264 400
rect 28896 0 28952 400
rect 33936 0 33992 400
<< obsm2 >>
rect 630 430 51674 52631
rect 630 400 25842 430
rect 25958 400 26178 430
rect 26294 400 28866 430
rect 28982 400 33906 430
rect 34022 400 51674 430
<< metal3 >>
rect 0 51744 400 51800
<< obsm3 >>
rect 400 51830 51679 52542
rect 430 51714 51679 51830
rect 400 1554 51679 51714
<< metal4 >>
rect 2224 1538 2384 52558
rect 9904 1538 10064 52558
rect 17584 1538 17744 52558
rect 25264 1538 25424 52558
rect 32944 1538 33104 52558
rect 40624 1538 40784 52558
rect 48304 1538 48464 52558
<< obsm4 >>
rect 1694 2193 2194 47759
rect 2414 2193 9874 47759
rect 10094 2193 17554 47759
rect 17774 2193 25234 47759
rect 25454 2193 32914 47759
rect 33134 2193 40594 47759
rect 40814 2193 48274 47759
rect 48494 2193 48706 47759
<< labels >>
rlabel metal2 s 25872 0 25928 400 6 spi_clock_i
port 1 nsew signal input
rlabel metal2 s 26208 0 26264 400 6 spi_cs_i
port 2 nsew signal input
rlabel metal2 s 33936 0 33992 400 6 spi_pico_i
port 3 nsew signal input
rlabel metal2 s 28896 0 28952 400 6 spi_poci_o
port 4 nsew signal output
rlabel metal3 s 0 51744 400 51800 6 sys_clock_i
port 5 nsew signal input
rlabel metal4 s 2224 1538 2384 52558 6 vdd
port 6 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 52558 6 vdd
port 6 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 52558 6 vdd
port 6 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 52558 6 vdd
port 6 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 52558 6 vss
port 7 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 52558 6 vss
port 7 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 52558 6 vss
port 7 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 52627 54419
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8633264
string GDS_FILE /home/kris/repos/diy-ic/lincoln-gfmpw-1d/openlane/titan/runs/23_12_08_11_53/results/signoff/titan.magic.gds
string GDS_START 410268
<< end >>

