magic
tech gf180mcuD
magscale 1 10
timestamp 1701901573
<< metal1 >>
rect 8754 38558 8766 38610
rect 8818 38607 8830 38610
rect 9762 38607 9774 38610
rect 8818 38561 9774 38607
rect 8818 38558 8830 38561
rect 9762 38558 9774 38561
rect 9826 38558 9838 38610
rect 12114 38558 12126 38610
rect 12178 38607 12190 38610
rect 13122 38607 13134 38610
rect 12178 38561 13134 38607
rect 12178 38558 12190 38561
rect 13122 38558 13134 38561
rect 13186 38558 13198 38610
rect 15922 38558 15934 38610
rect 15986 38607 15998 38610
rect 16706 38607 16718 38610
rect 15986 38561 16718 38607
rect 15986 38558 15998 38561
rect 16706 38558 16718 38561
rect 16770 38558 16782 38610
rect 25554 38558 25566 38610
rect 25618 38607 25630 38610
rect 26338 38607 26350 38610
rect 25618 38561 26350 38607
rect 25618 38558 25630 38561
rect 26338 38558 26350 38561
rect 26402 38558 26414 38610
rect 27010 38558 27022 38610
rect 27074 38607 27086 38610
rect 28466 38607 28478 38610
rect 27074 38561 28478 38607
rect 27074 38558 27086 38561
rect 28466 38558 28478 38561
rect 28530 38558 28542 38610
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 13134 38274 13186 38286
rect 13134 38210 13186 38222
rect 15486 38274 15538 38286
rect 15486 38210 15538 38222
rect 18174 38274 18226 38286
rect 18174 38210 18226 38222
rect 20190 38274 20242 38286
rect 20190 38210 20242 38222
rect 12686 38162 12738 38174
rect 9762 38110 9774 38162
rect 9826 38110 9838 38162
rect 12686 38098 12738 38110
rect 18734 38162 18786 38174
rect 21298 38110 21310 38162
rect 21362 38110 21374 38162
rect 22866 38110 22878 38162
rect 22930 38110 22942 38162
rect 24770 38110 24782 38162
rect 24834 38110 24846 38162
rect 26338 38110 26350 38162
rect 26402 38110 26414 38162
rect 28802 38110 28814 38162
rect 28866 38110 28878 38162
rect 30370 38110 30382 38162
rect 30434 38110 30446 38162
rect 32722 38110 32734 38162
rect 32786 38110 32798 38162
rect 34402 38110 34414 38162
rect 34466 38110 34478 38162
rect 18734 38098 18786 38110
rect 11006 38050 11058 38062
rect 11006 37986 11058 37998
rect 11678 38050 11730 38062
rect 17490 37998 17502 38050
rect 17554 37998 17566 38050
rect 22082 37998 22094 38050
rect 22146 37998 22158 38050
rect 23426 37998 23438 38050
rect 23490 37998 23502 38050
rect 25554 37998 25566 38050
rect 25618 37998 25630 38050
rect 27234 37998 27246 38050
rect 27298 37998 27310 38050
rect 28466 37998 28478 38050
rect 28530 37998 28542 38050
rect 33730 37998 33742 38050
rect 33794 37998 33806 38050
rect 35410 37998 35422 38050
rect 35474 37998 35486 38050
rect 11678 37986 11730 37998
rect 9326 37826 9378 37838
rect 9326 37762 9378 37774
rect 11454 37826 11506 37838
rect 13918 37826 13970 37838
rect 12002 37774 12014 37826
rect 12066 37774 12078 37826
rect 11454 37762 11506 37774
rect 13918 37762 13970 37774
rect 14814 37826 14866 37838
rect 14814 37762 14866 37774
rect 15262 37826 15314 37838
rect 15262 37762 15314 37774
rect 16270 37826 16322 37838
rect 16270 37762 16322 37774
rect 17166 37826 17218 37838
rect 17166 37762 17218 37774
rect 19182 37826 19234 37838
rect 19182 37762 19234 37774
rect 19406 37826 19458 37838
rect 19406 37762 19458 37774
rect 23998 37826 24050 37838
rect 23998 37762 24050 37774
rect 27806 37826 27858 37838
rect 27806 37762 27858 37774
rect 29710 37826 29762 37838
rect 29710 37762 29762 37774
rect 29934 37826 29986 37838
rect 29934 37762 29986 37774
rect 31278 37826 31330 37838
rect 31278 37762 31330 37774
rect 31614 37826 31666 37838
rect 31614 37762 31666 37774
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 9102 37490 9154 37502
rect 9102 37426 9154 37438
rect 9662 37490 9714 37502
rect 15934 37490 15986 37502
rect 14578 37438 14590 37490
rect 14642 37438 14654 37490
rect 9662 37426 9714 37438
rect 15934 37426 15986 37438
rect 17390 37490 17442 37502
rect 17390 37426 17442 37438
rect 18958 37490 19010 37502
rect 23214 37490 23266 37502
rect 22642 37438 22654 37490
rect 22706 37438 22718 37490
rect 18958 37426 19010 37438
rect 23214 37426 23266 37438
rect 23998 37490 24050 37502
rect 29598 37490 29650 37502
rect 28914 37438 28926 37490
rect 28978 37438 28990 37490
rect 23998 37426 24050 37438
rect 29598 37426 29650 37438
rect 32398 37490 32450 37502
rect 32398 37426 32450 37438
rect 34974 37490 35026 37502
rect 34974 37426 35026 37438
rect 25230 37378 25282 37390
rect 19282 37326 19294 37378
rect 19346 37326 19358 37378
rect 24322 37326 24334 37378
rect 24386 37326 24398 37378
rect 25230 37314 25282 37326
rect 25342 37378 25394 37390
rect 25342 37314 25394 37326
rect 31390 37378 31442 37390
rect 31390 37314 31442 37326
rect 11678 37266 11730 37278
rect 19518 37266 19570 37278
rect 24670 37266 24722 37278
rect 12114 37214 12126 37266
rect 12178 37214 12190 37266
rect 16706 37214 16718 37266
rect 16770 37214 16782 37266
rect 18050 37214 18062 37266
rect 18114 37214 18126 37266
rect 20178 37214 20190 37266
rect 20242 37214 20254 37266
rect 11678 37202 11730 37214
rect 19518 37202 19570 37214
rect 24670 37202 24722 37214
rect 25566 37266 25618 37278
rect 25566 37202 25618 37214
rect 25902 37266 25954 37278
rect 29822 37266 29874 37278
rect 31166 37266 31218 37278
rect 26562 37214 26574 37266
rect 26626 37214 26638 37266
rect 30258 37214 30270 37266
rect 30322 37214 30334 37266
rect 25902 37202 25954 37214
rect 29822 37202 29874 37214
rect 31166 37202 31218 37214
rect 31502 37266 31554 37278
rect 31502 37202 31554 37214
rect 33630 37266 33682 37278
rect 33630 37202 33682 37214
rect 10782 37154 10834 37166
rect 10098 37102 10110 37154
rect 10162 37102 10174 37154
rect 10782 37090 10834 37102
rect 11230 37154 11282 37166
rect 18622 37154 18674 37166
rect 15474 37102 15486 37154
rect 15538 37102 15550 37154
rect 16370 37102 16382 37154
rect 16434 37102 16446 37154
rect 11230 37090 11282 37102
rect 18622 37090 18674 37102
rect 23438 37154 23490 37166
rect 23438 37090 23490 37102
rect 30830 37154 30882 37166
rect 33294 37154 33346 37166
rect 31938 37102 31950 37154
rect 32002 37102 32014 37154
rect 30830 37090 30882 37102
rect 33294 37090 33346 37102
rect 34078 37154 34130 37166
rect 34078 37090 34130 37102
rect 34526 37154 34578 37166
rect 34526 37090 34578 37102
rect 15150 37042 15202 37054
rect 15150 36978 15202 36990
rect 30942 37042 30994 37054
rect 30942 36978 30994 36990
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 12574 36706 12626 36718
rect 12574 36642 12626 36654
rect 14926 36706 14978 36718
rect 14926 36642 14978 36654
rect 22878 36706 22930 36718
rect 22878 36642 22930 36654
rect 27246 36706 27298 36718
rect 27246 36642 27298 36654
rect 32734 36706 32786 36718
rect 32734 36642 32786 36654
rect 36542 36706 36594 36718
rect 36542 36642 36594 36654
rect 12910 36594 12962 36606
rect 12910 36530 12962 36542
rect 16158 36594 16210 36606
rect 16158 36530 16210 36542
rect 21422 36594 21474 36606
rect 21422 36530 21474 36542
rect 27582 36594 27634 36606
rect 27582 36530 27634 36542
rect 9102 36482 9154 36494
rect 16494 36482 16546 36494
rect 21982 36482 22034 36494
rect 9538 36430 9550 36482
rect 9602 36430 9614 36482
rect 15362 36430 15374 36482
rect 15426 36430 15438 36482
rect 17042 36430 17054 36482
rect 17106 36430 17118 36482
rect 9102 36418 9154 36430
rect 16494 36418 16546 36430
rect 21982 36418 22034 36430
rect 23550 36482 23602 36494
rect 28254 36482 28306 36494
rect 24210 36430 24222 36482
rect 24274 36430 24286 36482
rect 28018 36430 28030 36482
rect 28082 36430 28094 36482
rect 23550 36418 23602 36430
rect 28254 36418 28306 36430
rect 29038 36482 29090 36494
rect 32846 36482 32898 36494
rect 29698 36430 29710 36482
rect 29762 36430 29774 36482
rect 33394 36430 33406 36482
rect 33458 36430 33470 36482
rect 29038 36418 29090 36430
rect 32846 36418 32898 36430
rect 13470 36370 13522 36382
rect 13470 36306 13522 36318
rect 13806 36370 13858 36382
rect 13806 36306 13858 36318
rect 14590 36370 14642 36382
rect 20526 36370 20578 36382
rect 15698 36318 15710 36370
rect 15762 36318 15774 36370
rect 14590 36306 14642 36318
rect 20526 36306 20578 36318
rect 22990 36370 23042 36382
rect 22990 36306 23042 36318
rect 27470 36370 27522 36382
rect 27470 36306 27522 36318
rect 27694 36370 27746 36382
rect 27694 36306 27746 36318
rect 28478 36370 28530 36382
rect 28478 36306 28530 36318
rect 28590 36370 28642 36382
rect 28590 36306 28642 36318
rect 31950 36370 32002 36382
rect 31950 36306 32002 36318
rect 12798 36258 12850 36270
rect 11890 36206 11902 36258
rect 11954 36206 11966 36258
rect 12798 36194 12850 36206
rect 16270 36258 16322 36270
rect 20190 36258 20242 36270
rect 19618 36206 19630 36258
rect 19682 36206 19694 36258
rect 16270 36194 16322 36206
rect 20190 36194 20242 36206
rect 20414 36258 20466 36270
rect 20414 36194 20466 36206
rect 21310 36258 21362 36270
rect 21310 36194 21362 36206
rect 21534 36258 21586 36270
rect 21534 36194 21586 36206
rect 22206 36258 22258 36270
rect 22530 36206 22542 36258
rect 22594 36206 22606 36258
rect 26562 36206 26574 36258
rect 26626 36206 26638 36258
rect 35746 36206 35758 36258
rect 35810 36206 35822 36258
rect 22206 36194 22258 36206
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 11342 35922 11394 35934
rect 11342 35858 11394 35870
rect 12238 35922 12290 35934
rect 12238 35858 12290 35870
rect 13134 35922 13186 35934
rect 13134 35858 13186 35870
rect 13582 35922 13634 35934
rect 13582 35858 13634 35870
rect 14030 35922 14082 35934
rect 14030 35858 14082 35870
rect 21422 35922 21474 35934
rect 21422 35858 21474 35870
rect 21982 35922 22034 35934
rect 21982 35858 22034 35870
rect 22206 35922 22258 35934
rect 22206 35858 22258 35870
rect 22766 35922 22818 35934
rect 22766 35858 22818 35870
rect 25342 35922 25394 35934
rect 25342 35858 25394 35870
rect 25678 35922 25730 35934
rect 25678 35858 25730 35870
rect 26238 35922 26290 35934
rect 26238 35858 26290 35870
rect 26574 35922 26626 35934
rect 26574 35858 26626 35870
rect 28366 35922 28418 35934
rect 28366 35858 28418 35870
rect 28926 35922 28978 35934
rect 28926 35858 28978 35870
rect 29374 35922 29426 35934
rect 29374 35858 29426 35870
rect 29822 35922 29874 35934
rect 29822 35858 29874 35870
rect 30718 35922 30770 35934
rect 30718 35858 30770 35870
rect 30830 35922 30882 35934
rect 30830 35858 30882 35870
rect 31950 35922 32002 35934
rect 31950 35858 32002 35870
rect 33182 35922 33234 35934
rect 33182 35858 33234 35870
rect 34414 35922 34466 35934
rect 34414 35858 34466 35870
rect 12014 35810 12066 35822
rect 12014 35746 12066 35758
rect 13918 35810 13970 35822
rect 13918 35746 13970 35758
rect 14478 35810 14530 35822
rect 14478 35746 14530 35758
rect 14926 35810 14978 35822
rect 14926 35746 14978 35758
rect 15150 35810 15202 35822
rect 15150 35746 15202 35758
rect 15710 35810 15762 35822
rect 15710 35746 15762 35758
rect 15934 35810 15986 35822
rect 15934 35746 15986 35758
rect 16382 35810 16434 35822
rect 16382 35746 16434 35758
rect 19630 35810 19682 35822
rect 19630 35746 19682 35758
rect 23550 35810 23602 35822
rect 23550 35746 23602 35758
rect 23662 35810 23714 35822
rect 23662 35746 23714 35758
rect 24670 35810 24722 35822
rect 24670 35746 24722 35758
rect 27134 35810 27186 35822
rect 27134 35746 27186 35758
rect 11006 35698 11058 35710
rect 11006 35634 11058 35646
rect 11230 35698 11282 35710
rect 11230 35634 11282 35646
rect 11454 35698 11506 35710
rect 11454 35634 11506 35646
rect 11902 35698 11954 35710
rect 11902 35634 11954 35646
rect 12350 35698 12402 35710
rect 12350 35634 12402 35646
rect 14366 35698 14418 35710
rect 14366 35634 14418 35646
rect 14702 35698 14754 35710
rect 14702 35634 14754 35646
rect 16270 35698 16322 35710
rect 16270 35634 16322 35646
rect 16494 35698 16546 35710
rect 16494 35634 16546 35646
rect 16942 35698 16994 35710
rect 19742 35698 19794 35710
rect 21310 35698 21362 35710
rect 17826 35646 17838 35698
rect 17890 35646 17902 35698
rect 19170 35646 19182 35698
rect 19234 35646 19246 35698
rect 21074 35646 21086 35698
rect 21138 35646 21150 35698
rect 16942 35634 16994 35646
rect 19742 35634 19794 35646
rect 21310 35634 21362 35646
rect 21534 35698 21586 35710
rect 22318 35698 22370 35710
rect 21746 35646 21758 35698
rect 21810 35646 21822 35698
rect 21534 35634 21586 35646
rect 22318 35634 22370 35646
rect 22654 35698 22706 35710
rect 22654 35634 22706 35646
rect 23886 35698 23938 35710
rect 23886 35634 23938 35646
rect 24222 35698 24274 35710
rect 24222 35634 24274 35646
rect 25230 35698 25282 35710
rect 25230 35634 25282 35646
rect 25454 35698 25506 35710
rect 25454 35634 25506 35646
rect 26686 35698 26738 35710
rect 30606 35698 30658 35710
rect 31838 35698 31890 35710
rect 27346 35646 27358 35698
rect 27410 35646 27422 35698
rect 31154 35646 31166 35698
rect 31218 35646 31230 35698
rect 26686 35634 26738 35646
rect 30606 35634 30658 35646
rect 31838 35634 31890 35646
rect 32062 35698 32114 35710
rect 32062 35634 32114 35646
rect 32510 35698 32562 35710
rect 32510 35634 32562 35646
rect 32958 35698 33010 35710
rect 32958 35634 33010 35646
rect 33294 35698 33346 35710
rect 33294 35634 33346 35646
rect 33742 35698 33794 35710
rect 33742 35634 33794 35646
rect 9998 35586 10050 35598
rect 9998 35522 10050 35534
rect 10558 35586 10610 35598
rect 17390 35586 17442 35598
rect 18734 35586 18786 35598
rect 15138 35534 15150 35586
rect 15202 35534 15214 35586
rect 15698 35534 15710 35586
rect 15762 35534 15774 35586
rect 18162 35534 18174 35586
rect 18226 35534 18238 35586
rect 10558 35522 10610 35534
rect 17390 35522 17442 35534
rect 18734 35522 18786 35534
rect 20302 35586 20354 35598
rect 20302 35522 20354 35534
rect 20750 35586 20802 35598
rect 20750 35522 20802 35534
rect 27918 35586 27970 35598
rect 27918 35522 27970 35534
rect 28814 35586 28866 35598
rect 28814 35522 28866 35534
rect 30270 35586 30322 35598
rect 30270 35522 30322 35534
rect 34302 35586 34354 35598
rect 34302 35522 34354 35534
rect 34862 35586 34914 35598
rect 34862 35522 34914 35534
rect 22766 35474 22818 35486
rect 24558 35474 24610 35486
rect 23986 35422 23998 35474
rect 24050 35471 24062 35474
rect 24322 35471 24334 35474
rect 24050 35425 24334 35471
rect 24050 35422 24062 35425
rect 24322 35422 24334 35425
rect 24386 35422 24398 35474
rect 22766 35410 22818 35422
rect 24558 35410 24610 35422
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 15486 35138 15538 35150
rect 7298 35086 7310 35138
rect 7362 35135 7374 35138
rect 7970 35135 7982 35138
rect 7362 35089 7982 35135
rect 7362 35086 7374 35089
rect 7970 35086 7982 35089
rect 8034 35086 8046 35138
rect 15486 35074 15538 35086
rect 20750 35138 20802 35150
rect 25442 35086 25454 35138
rect 25506 35135 25518 35138
rect 26114 35135 26126 35138
rect 25506 35089 26126 35135
rect 25506 35086 25518 35089
rect 26114 35086 26126 35089
rect 26178 35086 26190 35138
rect 20750 35074 20802 35086
rect 7534 35026 7586 35038
rect 7534 34962 7586 34974
rect 7982 35026 8034 35038
rect 7982 34962 8034 34974
rect 8654 35026 8706 35038
rect 12462 35026 12514 35038
rect 19406 35026 19458 35038
rect 10546 34974 10558 35026
rect 10610 34974 10622 35026
rect 14802 34974 14814 35026
rect 14866 34974 14878 35026
rect 16258 34974 16270 35026
rect 16322 34974 16334 35026
rect 8654 34962 8706 34974
rect 12462 34962 12514 34974
rect 19406 34962 19458 34974
rect 19854 35026 19906 35038
rect 19854 34962 19906 34974
rect 20414 35026 20466 35038
rect 20414 34962 20466 34974
rect 20638 35026 20690 35038
rect 20638 34962 20690 34974
rect 22990 35026 23042 35038
rect 29710 35026 29762 35038
rect 24546 34974 24558 35026
rect 24610 34974 24622 35026
rect 22990 34962 23042 34974
rect 29710 34962 29762 34974
rect 30270 35026 30322 35038
rect 32510 35026 32562 35038
rect 31826 34974 31838 35026
rect 31890 34974 31902 35026
rect 30270 34962 30322 34974
rect 32510 34962 32562 34974
rect 33406 35026 33458 35038
rect 33406 34962 33458 34974
rect 7086 34914 7138 34926
rect 7086 34850 7138 34862
rect 8766 34914 8818 34926
rect 8766 34850 8818 34862
rect 9774 34914 9826 34926
rect 11902 34914 11954 34926
rect 10658 34862 10670 34914
rect 10722 34862 10734 34914
rect 11666 34862 11678 34914
rect 11730 34862 11742 34914
rect 9774 34850 9826 34862
rect 11902 34850 11954 34862
rect 14030 34914 14082 34926
rect 14030 34850 14082 34862
rect 14478 34914 14530 34926
rect 14478 34850 14530 34862
rect 16046 34914 16098 34926
rect 16830 34914 16882 34926
rect 17726 34914 17778 34926
rect 16482 34862 16494 34914
rect 16546 34862 16558 34914
rect 17490 34862 17502 34914
rect 17554 34862 17566 34914
rect 16046 34850 16098 34862
rect 16830 34850 16882 34862
rect 17726 34850 17778 34862
rect 18062 34914 18114 34926
rect 18062 34850 18114 34862
rect 18398 34914 18450 34926
rect 23214 34914 23266 34926
rect 22194 34862 22206 34914
rect 22258 34862 22270 34914
rect 22418 34862 22430 34914
rect 22482 34862 22494 34914
rect 18398 34850 18450 34862
rect 23214 34850 23266 34862
rect 23438 34914 23490 34926
rect 23438 34850 23490 34862
rect 24222 34914 24274 34926
rect 24222 34850 24274 34862
rect 25678 34914 25730 34926
rect 25678 34850 25730 34862
rect 27134 34914 27186 34926
rect 33966 34914 34018 34926
rect 31378 34862 31390 34914
rect 31442 34862 31454 34914
rect 32050 34862 32062 34914
rect 32114 34862 32126 34914
rect 27134 34850 27186 34862
rect 33966 34850 34018 34862
rect 9998 34802 10050 34814
rect 9998 34738 10050 34750
rect 11006 34802 11058 34814
rect 11006 34738 11058 34750
rect 13918 34802 13970 34814
rect 13918 34738 13970 34750
rect 14142 34802 14194 34814
rect 14142 34738 14194 34750
rect 15822 34802 15874 34814
rect 15822 34738 15874 34750
rect 18286 34802 18338 34814
rect 18286 34738 18338 34750
rect 18846 34802 18898 34814
rect 18846 34738 18898 34750
rect 18958 34802 19010 34814
rect 18958 34738 19010 34750
rect 22654 34802 22706 34814
rect 22654 34738 22706 34750
rect 24558 34802 24610 34814
rect 24558 34738 24610 34750
rect 25230 34802 25282 34814
rect 25230 34738 25282 34750
rect 26574 34802 26626 34814
rect 26574 34738 26626 34750
rect 26910 34802 26962 34814
rect 26910 34738 26962 34750
rect 28142 34802 28194 34814
rect 28142 34738 28194 34750
rect 28254 34802 28306 34814
rect 28254 34738 28306 34750
rect 32398 34802 32450 34814
rect 32398 34738 32450 34750
rect 32734 34802 32786 34814
rect 32734 34738 32786 34750
rect 32958 34802 33010 34814
rect 32958 34738 33010 34750
rect 6750 34690 6802 34702
rect 6750 34626 6802 34638
rect 6974 34690 7026 34702
rect 6974 34626 7026 34638
rect 9102 34690 9154 34702
rect 9102 34626 9154 34638
rect 9214 34690 9266 34702
rect 9214 34626 9266 34638
rect 9326 34690 9378 34702
rect 9326 34626 9378 34638
rect 10222 34690 10274 34702
rect 10222 34626 10274 34638
rect 10446 34690 10498 34702
rect 10446 34626 10498 34638
rect 13022 34690 13074 34702
rect 13022 34626 13074 34638
rect 14702 34690 14754 34702
rect 14702 34626 14754 34638
rect 15262 34690 15314 34702
rect 15262 34626 15314 34638
rect 15374 34690 15426 34702
rect 15374 34626 15426 34638
rect 16270 34690 16322 34702
rect 16270 34626 16322 34638
rect 18622 34690 18674 34702
rect 18622 34626 18674 34638
rect 23886 34690 23938 34702
rect 23886 34626 23938 34638
rect 24334 34690 24386 34702
rect 24334 34626 24386 34638
rect 24670 34690 24722 34702
rect 24670 34626 24722 34638
rect 26126 34690 26178 34702
rect 26126 34626 26178 34638
rect 27246 34690 27298 34702
rect 27246 34626 27298 34638
rect 27358 34690 27410 34702
rect 27358 34626 27410 34638
rect 27470 34690 27522 34702
rect 27470 34626 27522 34638
rect 27918 34690 27970 34702
rect 27918 34626 27970 34638
rect 29374 34690 29426 34702
rect 29374 34626 29426 34638
rect 30942 34690 30994 34702
rect 30942 34626 30994 34638
rect 31614 34690 31666 34702
rect 31614 34626 31666 34638
rect 31838 34690 31890 34702
rect 31838 34626 31890 34638
rect 33518 34690 33570 34702
rect 33518 34626 33570 34638
rect 34414 34690 34466 34702
rect 34414 34626 34466 34638
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 7422 34354 7474 34366
rect 7422 34290 7474 34302
rect 14478 34354 14530 34366
rect 14478 34290 14530 34302
rect 14702 34354 14754 34366
rect 14702 34290 14754 34302
rect 14926 34354 14978 34366
rect 14926 34290 14978 34302
rect 16942 34354 16994 34366
rect 16942 34290 16994 34302
rect 17502 34354 17554 34366
rect 17502 34290 17554 34302
rect 18510 34354 18562 34366
rect 18510 34290 18562 34302
rect 18734 34354 18786 34366
rect 18734 34290 18786 34302
rect 25454 34354 25506 34366
rect 25454 34290 25506 34302
rect 29374 34354 29426 34366
rect 29374 34290 29426 34302
rect 30718 34354 30770 34366
rect 30718 34290 30770 34302
rect 30830 34354 30882 34366
rect 30830 34290 30882 34302
rect 6638 34242 6690 34254
rect 6638 34178 6690 34190
rect 11342 34242 11394 34254
rect 11342 34178 11394 34190
rect 13918 34242 13970 34254
rect 13918 34178 13970 34190
rect 16718 34242 16770 34254
rect 16718 34178 16770 34190
rect 21086 34242 21138 34254
rect 21086 34178 21138 34190
rect 21422 34242 21474 34254
rect 21422 34178 21474 34190
rect 25678 34242 25730 34254
rect 25678 34178 25730 34190
rect 27582 34242 27634 34254
rect 27582 34178 27634 34190
rect 27918 34242 27970 34254
rect 27918 34178 27970 34190
rect 31390 34242 31442 34254
rect 31390 34178 31442 34190
rect 3950 34130 4002 34142
rect 8878 34130 8930 34142
rect 4274 34078 4286 34130
rect 4338 34078 4350 34130
rect 8530 34078 8542 34130
rect 8594 34078 8606 34130
rect 3950 34066 4002 34078
rect 8878 34066 8930 34078
rect 10110 34130 10162 34142
rect 11454 34130 11506 34142
rect 14030 34130 14082 34142
rect 10770 34078 10782 34130
rect 10834 34078 10846 34130
rect 12002 34078 12014 34130
rect 12066 34078 12078 34130
rect 12674 34078 12686 34130
rect 12738 34078 12750 34130
rect 10110 34066 10162 34078
rect 11454 34066 11506 34078
rect 14030 34066 14082 34078
rect 15374 34130 15426 34142
rect 16606 34130 16658 34142
rect 15586 34078 15598 34130
rect 15650 34078 15662 34130
rect 15374 34066 15426 34078
rect 16606 34066 16658 34078
rect 17390 34130 17442 34142
rect 19182 34130 19234 34142
rect 20974 34130 21026 34142
rect 22318 34130 22370 34142
rect 24110 34130 24162 34142
rect 17602 34078 17614 34130
rect 17666 34078 17678 34130
rect 20626 34078 20638 34130
rect 20690 34078 20702 34130
rect 22082 34078 22094 34130
rect 22146 34078 22158 34130
rect 23314 34078 23326 34130
rect 23378 34078 23390 34130
rect 17390 34066 17442 34078
rect 19182 34066 19234 34078
rect 20974 34066 21026 34078
rect 22318 34066 22370 34078
rect 24110 34066 24162 34078
rect 24334 34130 24386 34142
rect 25230 34130 25282 34142
rect 24658 34078 24670 34130
rect 24722 34078 24734 34130
rect 24334 34066 24386 34078
rect 25230 34066 25282 34078
rect 26238 34130 26290 34142
rect 28030 34130 28082 34142
rect 30494 34130 30546 34142
rect 27122 34078 27134 34130
rect 27186 34078 27198 34130
rect 27346 34078 27358 34130
rect 27410 34078 27422 34130
rect 28466 34078 28478 34130
rect 28530 34078 28542 34130
rect 26238 34066 26290 34078
rect 28030 34066 28082 34078
rect 30494 34066 30546 34078
rect 30606 34130 30658 34142
rect 31042 34078 31054 34130
rect 31106 34078 31118 34130
rect 32274 34078 32286 34130
rect 32338 34078 32350 34130
rect 33618 34078 33630 34130
rect 33682 34078 33694 34130
rect 30606 34066 30658 34078
rect 8990 34018 9042 34030
rect 14814 34018 14866 34030
rect 12786 33966 12798 34018
rect 12850 33966 12862 34018
rect 8990 33954 9042 33966
rect 14814 33954 14866 33966
rect 16270 34018 16322 34030
rect 16270 33954 16322 33966
rect 18622 34018 18674 34030
rect 18622 33954 18674 33966
rect 19518 34018 19570 34030
rect 23774 34018 23826 34030
rect 23426 33966 23438 34018
rect 23490 33966 23502 34018
rect 19518 33954 19570 33966
rect 23774 33954 23826 33966
rect 24222 34018 24274 34030
rect 24222 33954 24274 33966
rect 25342 34018 25394 34030
rect 25342 33954 25394 33966
rect 26126 34018 26178 34030
rect 26126 33954 26178 33966
rect 29822 34018 29874 34030
rect 34078 34018 34130 34030
rect 32162 33966 32174 34018
rect 32226 33966 32238 34018
rect 33282 33966 33294 34018
rect 33346 33966 33358 34018
rect 29822 33954 29874 33966
rect 34078 33954 34130 33966
rect 13918 33906 13970 33918
rect 10210 33854 10222 33906
rect 10274 33854 10286 33906
rect 13918 33842 13970 33854
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 6974 33570 7026 33582
rect 6974 33506 7026 33518
rect 10558 33570 10610 33582
rect 14590 33570 14642 33582
rect 27918 33570 27970 33582
rect 12114 33518 12126 33570
rect 12178 33518 12190 33570
rect 24546 33518 24558 33570
rect 24610 33518 24622 33570
rect 10558 33506 10610 33518
rect 14590 33506 14642 33518
rect 27918 33506 27970 33518
rect 6190 33458 6242 33470
rect 6190 33394 6242 33406
rect 8094 33458 8146 33470
rect 8094 33394 8146 33406
rect 9998 33458 10050 33470
rect 9998 33394 10050 33406
rect 15038 33458 15090 33470
rect 16494 33458 16546 33470
rect 15810 33406 15822 33458
rect 15874 33406 15886 33458
rect 15038 33394 15090 33406
rect 16494 33394 16546 33406
rect 19070 33458 19122 33470
rect 19070 33394 19122 33406
rect 23662 33458 23714 33470
rect 23662 33394 23714 33406
rect 26126 33458 26178 33470
rect 27582 33458 27634 33470
rect 31950 33458 32002 33470
rect 27122 33406 27134 33458
rect 27186 33406 27198 33458
rect 28242 33406 28254 33458
rect 28306 33406 28318 33458
rect 31602 33406 31614 33458
rect 31666 33406 31678 33458
rect 26126 33394 26178 33406
rect 27582 33394 27634 33406
rect 31950 33394 32002 33406
rect 33630 33458 33682 33470
rect 33630 33394 33682 33406
rect 7870 33346 7922 33358
rect 6626 33294 6638 33346
rect 6690 33294 6702 33346
rect 7870 33282 7922 33294
rect 8878 33346 8930 33358
rect 10894 33346 10946 33358
rect 9650 33294 9662 33346
rect 9714 33294 9726 33346
rect 8878 33282 8930 33294
rect 10894 33282 10946 33294
rect 11454 33346 11506 33358
rect 14702 33346 14754 33358
rect 16382 33346 16434 33358
rect 11666 33294 11678 33346
rect 11730 33294 11742 33346
rect 15474 33294 15486 33346
rect 15538 33294 15550 33346
rect 11454 33282 11506 33294
rect 14702 33282 14754 33294
rect 16382 33282 16434 33294
rect 16606 33346 16658 33358
rect 16606 33282 16658 33294
rect 17054 33346 17106 33358
rect 18846 33346 18898 33358
rect 17602 33294 17614 33346
rect 17666 33294 17678 33346
rect 17054 33282 17106 33294
rect 18846 33282 18898 33294
rect 21758 33346 21810 33358
rect 21758 33282 21810 33294
rect 21982 33346 22034 33358
rect 21982 33282 22034 33294
rect 22430 33346 22482 33358
rect 23550 33346 23602 33358
rect 23202 33294 23214 33346
rect 23266 33294 23278 33346
rect 22430 33282 22482 33294
rect 23550 33282 23602 33294
rect 23998 33346 24050 33358
rect 23998 33282 24050 33294
rect 24222 33346 24274 33358
rect 24222 33282 24274 33294
rect 25118 33346 25170 33358
rect 30382 33346 30434 33358
rect 33182 33346 33234 33358
rect 26898 33294 26910 33346
rect 26962 33294 26974 33346
rect 31490 33294 31502 33346
rect 31554 33294 31566 33346
rect 32722 33294 32734 33346
rect 32786 33294 32798 33346
rect 25118 33282 25170 33294
rect 30382 33282 30434 33294
rect 33182 33282 33234 33294
rect 33742 33346 33794 33358
rect 35086 33346 35138 33358
rect 34178 33294 34190 33346
rect 34242 33294 34254 33346
rect 35298 33294 35310 33346
rect 35362 33294 35374 33346
rect 33742 33282 33794 33294
rect 35086 33282 35138 33294
rect 7086 33234 7138 33246
rect 7086 33170 7138 33182
rect 8542 33234 8594 33246
rect 8542 33170 8594 33182
rect 9102 33234 9154 33246
rect 9102 33170 9154 33182
rect 11118 33234 11170 33246
rect 18734 33234 18786 33246
rect 17826 33182 17838 33234
rect 17890 33182 17902 33234
rect 18386 33182 18398 33234
rect 18450 33182 18462 33234
rect 11118 33170 11170 33182
rect 18734 33170 18786 33182
rect 21870 33234 21922 33246
rect 21870 33170 21922 33182
rect 25006 33234 25058 33246
rect 25006 33170 25058 33182
rect 28142 33234 28194 33246
rect 28142 33170 28194 33182
rect 30494 33234 30546 33246
rect 30494 33170 30546 33182
rect 32286 33234 32338 33246
rect 32286 33170 32338 33182
rect 34974 33234 35026 33246
rect 34974 33170 35026 33182
rect 6078 33122 6130 33134
rect 6078 33058 6130 33070
rect 6302 33122 6354 33134
rect 6302 33058 6354 33070
rect 8206 33122 8258 33134
rect 8206 33058 8258 33070
rect 8654 33122 8706 33134
rect 8654 33058 8706 33070
rect 9550 33122 9602 33134
rect 9550 33058 9602 33070
rect 19182 33122 19234 33134
rect 19182 33058 19234 33070
rect 19406 33122 19458 33134
rect 19406 33058 19458 33070
rect 19966 33122 20018 33134
rect 19966 33058 20018 33070
rect 24782 33122 24834 33134
rect 24782 33058 24834 33070
rect 26238 33122 26290 33134
rect 26238 33058 26290 33070
rect 30718 33122 30770 33134
rect 30718 33058 30770 33070
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 13582 32786 13634 32798
rect 13582 32722 13634 32734
rect 15150 32786 15202 32798
rect 15150 32722 15202 32734
rect 16830 32786 16882 32798
rect 16830 32722 16882 32734
rect 23326 32786 23378 32798
rect 23326 32722 23378 32734
rect 27134 32786 27186 32798
rect 27134 32722 27186 32734
rect 30830 32786 30882 32798
rect 30830 32722 30882 32734
rect 33406 32786 33458 32798
rect 33406 32722 33458 32734
rect 8654 32674 8706 32686
rect 8654 32610 8706 32622
rect 9998 32674 10050 32686
rect 9998 32610 10050 32622
rect 10446 32674 10498 32686
rect 10446 32610 10498 32622
rect 10894 32674 10946 32686
rect 10894 32610 10946 32622
rect 12574 32674 12626 32686
rect 12574 32610 12626 32622
rect 13694 32674 13746 32686
rect 22654 32674 22706 32686
rect 18274 32622 18286 32674
rect 18338 32622 18350 32674
rect 19282 32622 19294 32674
rect 19346 32622 19358 32674
rect 13694 32610 13746 32622
rect 22654 32610 22706 32622
rect 24110 32674 24162 32686
rect 24110 32610 24162 32622
rect 26910 32674 26962 32686
rect 26910 32610 26962 32622
rect 27918 32674 27970 32686
rect 27918 32610 27970 32622
rect 28030 32674 28082 32686
rect 28030 32610 28082 32622
rect 30606 32674 30658 32686
rect 30606 32610 30658 32622
rect 31054 32674 31106 32686
rect 31054 32610 31106 32622
rect 34078 32674 34130 32686
rect 34078 32610 34130 32622
rect 9886 32562 9938 32574
rect 8194 32510 8206 32562
rect 8258 32510 8270 32562
rect 9886 32498 9938 32510
rect 10110 32562 10162 32574
rect 10110 32498 10162 32510
rect 10670 32562 10722 32574
rect 10670 32498 10722 32510
rect 11006 32562 11058 32574
rect 11006 32498 11058 32510
rect 12798 32562 12850 32574
rect 12798 32498 12850 32510
rect 14702 32562 14754 32574
rect 14702 32498 14754 32510
rect 14926 32562 14978 32574
rect 22766 32562 22818 32574
rect 17714 32510 17726 32562
rect 17778 32510 17790 32562
rect 19394 32510 19406 32562
rect 19458 32510 19470 32562
rect 14926 32498 14978 32510
rect 22766 32498 22818 32510
rect 23214 32562 23266 32574
rect 23214 32498 23266 32510
rect 23550 32562 23602 32574
rect 23550 32498 23602 32510
rect 23998 32562 24050 32574
rect 23998 32498 24050 32510
rect 24222 32562 24274 32574
rect 24222 32498 24274 32510
rect 24670 32562 24722 32574
rect 24670 32498 24722 32510
rect 27246 32562 27298 32574
rect 27246 32498 27298 32510
rect 27358 32562 27410 32574
rect 27358 32498 27410 32510
rect 30494 32562 30546 32574
rect 32958 32562 33010 32574
rect 31714 32510 31726 32562
rect 31778 32510 31790 32562
rect 30494 32498 30546 32510
rect 32958 32498 33010 32510
rect 33630 32562 33682 32574
rect 33630 32498 33682 32510
rect 33854 32562 33906 32574
rect 33854 32498 33906 32510
rect 34190 32562 34242 32574
rect 34190 32498 34242 32510
rect 6078 32450 6130 32462
rect 6078 32386 6130 32398
rect 6862 32450 6914 32462
rect 6862 32386 6914 32398
rect 7310 32450 7362 32462
rect 11454 32450 11506 32462
rect 7746 32398 7758 32450
rect 7810 32398 7822 32450
rect 7310 32386 7362 32398
rect 11454 32386 11506 32398
rect 14142 32450 14194 32462
rect 14142 32386 14194 32398
rect 14814 32450 14866 32462
rect 14814 32386 14866 32398
rect 16382 32450 16434 32462
rect 33518 32450 33570 32462
rect 20962 32398 20974 32450
rect 21026 32398 21038 32450
rect 31378 32398 31390 32450
rect 31442 32398 31454 32450
rect 16382 32386 16434 32398
rect 33518 32386 33570 32398
rect 13134 32338 13186 32350
rect 13134 32274 13186 32286
rect 13582 32338 13634 32350
rect 13582 32274 13634 32286
rect 14030 32338 14082 32350
rect 14030 32274 14082 32286
rect 27918 32338 27970 32350
rect 27918 32274 27970 32286
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 7758 32002 7810 32014
rect 7758 31938 7810 31950
rect 5854 31890 5906 31902
rect 5854 31826 5906 31838
rect 6302 31890 6354 31902
rect 6302 31826 6354 31838
rect 6862 31890 6914 31902
rect 6862 31826 6914 31838
rect 19406 31890 19458 31902
rect 19406 31826 19458 31838
rect 24222 31890 24274 31902
rect 24222 31826 24274 31838
rect 26350 31890 26402 31902
rect 26350 31826 26402 31838
rect 28030 31890 28082 31902
rect 28030 31826 28082 31838
rect 28478 31890 28530 31902
rect 30930 31838 30942 31890
rect 30994 31838 31006 31890
rect 33170 31838 33182 31890
rect 33234 31838 33246 31890
rect 28478 31826 28530 31838
rect 18622 31778 18674 31790
rect 22430 31778 22482 31790
rect 7746 31726 7758 31778
rect 7810 31726 7822 31778
rect 13570 31726 13582 31778
rect 13634 31726 13646 31778
rect 15250 31726 15262 31778
rect 15314 31726 15326 31778
rect 17266 31726 17278 31778
rect 17330 31726 17342 31778
rect 22194 31726 22206 31778
rect 22258 31726 22270 31778
rect 18622 31714 18674 31726
rect 22430 31714 22482 31726
rect 23438 31778 23490 31790
rect 23438 31714 23490 31726
rect 23886 31778 23938 31790
rect 25678 31778 25730 31790
rect 24434 31726 24446 31778
rect 24498 31726 24510 31778
rect 23886 31714 23938 31726
rect 25678 31714 25730 31726
rect 26574 31778 26626 31790
rect 26574 31714 26626 31726
rect 27022 31778 27074 31790
rect 27022 31714 27074 31726
rect 27918 31778 27970 31790
rect 27918 31714 27970 31726
rect 28142 31778 28194 31790
rect 31278 31778 31330 31790
rect 29138 31726 29150 31778
rect 29202 31726 29214 31778
rect 28142 31714 28194 31726
rect 31278 31714 31330 31726
rect 31838 31778 31890 31790
rect 31838 31714 31890 31726
rect 32062 31778 32114 31790
rect 32062 31714 32114 31726
rect 32510 31778 32562 31790
rect 32510 31714 32562 31726
rect 33742 31778 33794 31790
rect 33742 31714 33794 31726
rect 7310 31666 7362 31678
rect 2034 31614 2046 31666
rect 2098 31614 2110 31666
rect 7310 31602 7362 31614
rect 8094 31666 8146 31678
rect 8094 31602 8146 31614
rect 8878 31666 8930 31678
rect 8878 31602 8930 31614
rect 9214 31666 9266 31678
rect 9214 31602 9266 31614
rect 11454 31666 11506 31678
rect 11454 31602 11506 31614
rect 11566 31666 11618 31678
rect 18398 31666 18450 31678
rect 13458 31614 13470 31666
rect 13522 31614 13534 31666
rect 15586 31614 15598 31666
rect 15650 31614 15662 31666
rect 17042 31614 17054 31666
rect 17106 31614 17118 31666
rect 11566 31602 11618 31614
rect 18398 31602 18450 31614
rect 19294 31666 19346 31678
rect 19294 31602 19346 31614
rect 23214 31666 23266 31678
rect 23214 31602 23266 31614
rect 24110 31666 24162 31678
rect 24110 31602 24162 31614
rect 26014 31666 26066 31678
rect 26014 31602 26066 31614
rect 26910 31666 26962 31678
rect 26910 31602 26962 31614
rect 27582 31666 27634 31678
rect 27582 31602 27634 31614
rect 28590 31666 28642 31678
rect 30606 31666 30658 31678
rect 29250 31614 29262 31666
rect 29314 31614 29326 31666
rect 29810 31614 29822 31666
rect 29874 31614 29886 31666
rect 28590 31602 28642 31614
rect 30606 31602 30658 31614
rect 30830 31666 30882 31678
rect 30830 31602 30882 31614
rect 31502 31666 31554 31678
rect 31502 31602 31554 31614
rect 32734 31666 32786 31678
rect 32734 31602 32786 31614
rect 33406 31666 33458 31678
rect 33406 31602 33458 31614
rect 33854 31666 33906 31678
rect 33854 31602 33906 31614
rect 39566 31666 39618 31678
rect 39566 31602 39618 31614
rect 1710 31554 1762 31566
rect 1710 31490 1762 31502
rect 2494 31554 2546 31566
rect 2494 31490 2546 31502
rect 5742 31554 5794 31566
rect 5742 31490 5794 31502
rect 7422 31554 7474 31566
rect 7422 31490 7474 31502
rect 8542 31554 8594 31566
rect 8542 31490 8594 31502
rect 8766 31554 8818 31566
rect 8766 31490 8818 31502
rect 9326 31554 9378 31566
rect 9326 31490 9378 31502
rect 9550 31554 9602 31566
rect 9550 31490 9602 31502
rect 11790 31554 11842 31566
rect 11790 31490 11842 31502
rect 18734 31554 18786 31566
rect 18734 31490 18786 31502
rect 18846 31554 18898 31566
rect 18846 31490 18898 31502
rect 22766 31554 22818 31566
rect 22766 31490 22818 31502
rect 23326 31554 23378 31566
rect 23326 31490 23378 31502
rect 25902 31554 25954 31566
rect 25902 31490 25954 31502
rect 26798 31554 26850 31566
rect 26798 31490 26850 31502
rect 31726 31554 31778 31566
rect 31726 31490 31778 31502
rect 32286 31554 32338 31566
rect 32286 31490 32338 31502
rect 34078 31554 34130 31566
rect 40238 31554 40290 31566
rect 39218 31502 39230 31554
rect 39282 31502 39294 31554
rect 39890 31502 39902 31554
rect 39954 31502 39966 31554
rect 34078 31490 34130 31502
rect 40238 31490 40290 31502
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 11118 31218 11170 31230
rect 3266 31166 3278 31218
rect 3330 31166 3342 31218
rect 10546 31166 10558 31218
rect 10610 31166 10622 31218
rect 11118 31154 11170 31166
rect 14702 31218 14754 31230
rect 14702 31154 14754 31166
rect 15374 31218 15426 31230
rect 15374 31154 15426 31166
rect 15598 31218 15650 31230
rect 15598 31154 15650 31166
rect 16718 31218 16770 31230
rect 16718 31154 16770 31166
rect 19518 31218 19570 31230
rect 19518 31154 19570 31166
rect 20750 31218 20802 31230
rect 20750 31154 20802 31166
rect 26126 31218 26178 31230
rect 26126 31154 26178 31166
rect 31614 31218 31666 31230
rect 31614 31154 31666 31166
rect 33070 31218 33122 31230
rect 33070 31154 33122 31166
rect 39902 31218 39954 31230
rect 39902 31154 39954 31166
rect 6526 31106 6578 31118
rect 6526 31042 6578 31054
rect 6638 31106 6690 31118
rect 6638 31042 6690 31054
rect 8542 31106 8594 31118
rect 8542 31042 8594 31054
rect 8766 31106 8818 31118
rect 8766 31042 8818 31054
rect 9550 31106 9602 31118
rect 16606 31106 16658 31118
rect 13458 31054 13470 31106
rect 13522 31054 13534 31106
rect 13794 31054 13806 31106
rect 13858 31054 13870 31106
rect 9550 31042 9602 31054
rect 16606 31042 16658 31054
rect 16830 31106 16882 31118
rect 16830 31042 16882 31054
rect 18510 31106 18562 31118
rect 18510 31042 18562 31054
rect 20638 31106 20690 31118
rect 20638 31042 20690 31054
rect 31502 31106 31554 31118
rect 31502 31042 31554 31054
rect 33294 31106 33346 31118
rect 33294 31042 33346 31054
rect 6190 30994 6242 31006
rect 8094 30994 8146 31006
rect 5618 30942 5630 30994
rect 5682 30942 5694 30994
rect 7746 30942 7758 30994
rect 7810 30942 7822 30994
rect 6190 30930 6242 30942
rect 8094 30930 8146 30942
rect 9662 30994 9714 31006
rect 9662 30930 9714 30942
rect 9886 30994 9938 31006
rect 9886 30930 9938 30942
rect 10110 30994 10162 31006
rect 10110 30930 10162 30942
rect 11006 30994 11058 31006
rect 11006 30930 11058 30942
rect 11342 30994 11394 31006
rect 11342 30930 11394 30942
rect 11454 30994 11506 31006
rect 15486 30994 15538 31006
rect 12114 30942 12126 30994
rect 12178 30942 12190 30994
rect 13010 30942 13022 30994
rect 13074 30942 13086 30994
rect 13906 30942 13918 30994
rect 13970 30942 13982 30994
rect 15026 30942 15038 30994
rect 15090 30942 15102 30994
rect 11454 30930 11506 30942
rect 15486 30930 15538 30942
rect 17502 30994 17554 31006
rect 17502 30930 17554 30942
rect 17950 30994 18002 31006
rect 17950 30930 18002 30942
rect 18174 30994 18226 31006
rect 18958 30994 19010 31006
rect 18722 30942 18734 30994
rect 18786 30942 18798 30994
rect 18174 30930 18226 30942
rect 18958 30930 19010 30942
rect 19406 30994 19458 31006
rect 19406 30930 19458 30942
rect 19966 30994 20018 31006
rect 22878 30994 22930 31006
rect 20962 30942 20974 30994
rect 21026 30942 21038 30994
rect 19966 30930 20018 30942
rect 22878 30930 22930 30942
rect 26014 30994 26066 31006
rect 32174 30994 32226 31006
rect 26786 30942 26798 30994
rect 26850 30942 26862 30994
rect 28466 30942 28478 30994
rect 28530 30942 28542 30994
rect 26014 30930 26066 30942
rect 32174 30930 32226 30942
rect 32398 30994 32450 31006
rect 32398 30930 32450 30942
rect 33742 30994 33794 31006
rect 33742 30930 33794 30942
rect 40238 30994 40290 31006
rect 40238 30930 40290 30942
rect 7198 30882 7250 30894
rect 14590 30882 14642 30894
rect 8866 30830 8878 30882
rect 8930 30830 8942 30882
rect 14242 30830 14254 30882
rect 14306 30830 14318 30882
rect 7198 30818 7250 30830
rect 14590 30818 14642 30830
rect 17726 30882 17778 30894
rect 17726 30818 17778 30830
rect 19182 30882 19234 30894
rect 19182 30818 19234 30830
rect 19742 30882 19794 30894
rect 19742 30818 19794 30830
rect 22542 30882 22594 30894
rect 27470 30882 27522 30894
rect 23314 30830 23326 30882
rect 23378 30830 23390 30882
rect 27010 30830 27022 30882
rect 27074 30830 27086 30882
rect 22542 30818 22594 30830
rect 27470 30818 27522 30830
rect 27806 30882 27858 30894
rect 30718 30882 30770 30894
rect 28242 30830 28254 30882
rect 28306 30830 28318 30882
rect 27806 30818 27858 30830
rect 30718 30818 30770 30830
rect 31278 30882 31330 30894
rect 31278 30818 31330 30830
rect 32062 30882 32114 30894
rect 32062 30818 32114 30830
rect 33182 30882 33234 30894
rect 33182 30818 33234 30830
rect 2494 30770 2546 30782
rect 2494 30706 2546 30718
rect 6526 30770 6578 30782
rect 32510 30770 32562 30782
rect 20290 30718 20302 30770
rect 20354 30718 20366 30770
rect 6526 30706 6578 30718
rect 32510 30706 32562 30718
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 14254 30434 14306 30446
rect 14254 30370 14306 30382
rect 18286 30434 18338 30446
rect 18286 30370 18338 30382
rect 21310 30434 21362 30446
rect 21310 30370 21362 30382
rect 26126 30434 26178 30446
rect 26126 30370 26178 30382
rect 10446 30322 10498 30334
rect 8082 30270 8094 30322
rect 8146 30270 8158 30322
rect 9762 30270 9774 30322
rect 9826 30270 9838 30322
rect 10446 30258 10498 30270
rect 14030 30322 14082 30334
rect 18174 30322 18226 30334
rect 21422 30322 21474 30334
rect 15362 30270 15374 30322
rect 15426 30270 15438 30322
rect 17378 30270 17390 30322
rect 17442 30270 17454 30322
rect 19394 30270 19406 30322
rect 19458 30270 19470 30322
rect 14030 30258 14082 30270
rect 18174 30258 18226 30270
rect 21422 30258 21474 30270
rect 2158 30210 2210 30222
rect 6078 30210 6130 30222
rect 2818 30158 2830 30210
rect 2882 30158 2894 30210
rect 2158 30146 2210 30158
rect 6078 30146 6130 30158
rect 6750 30210 6802 30222
rect 11902 30210 11954 30222
rect 6962 30158 6974 30210
rect 7026 30158 7038 30210
rect 8194 30158 8206 30210
rect 8258 30158 8270 30210
rect 8866 30158 8878 30210
rect 8930 30158 8942 30210
rect 9314 30158 9326 30210
rect 9378 30158 9390 30210
rect 10210 30158 10222 30210
rect 10274 30158 10286 30210
rect 6750 30146 6802 30158
rect 11902 30146 11954 30158
rect 12238 30210 12290 30222
rect 12238 30146 12290 30158
rect 12462 30210 12514 30222
rect 12462 30146 12514 30158
rect 12798 30210 12850 30222
rect 12798 30146 12850 30158
rect 13806 30210 13858 30222
rect 13806 30146 13858 30158
rect 14478 30210 14530 30222
rect 18622 30210 18674 30222
rect 20078 30210 20130 30222
rect 15474 30158 15486 30210
rect 15538 30158 15550 30210
rect 17154 30158 17166 30210
rect 17218 30158 17230 30210
rect 17938 30158 17950 30210
rect 18002 30158 18014 30210
rect 19170 30158 19182 30210
rect 19234 30158 19246 30210
rect 14478 30146 14530 30158
rect 18622 30146 18674 30158
rect 20078 30146 20130 30158
rect 20526 30210 20578 30222
rect 22766 30210 22818 30222
rect 27470 30210 27522 30222
rect 29150 30210 29202 30222
rect 21634 30158 21646 30210
rect 21698 30158 21710 30210
rect 23314 30158 23326 30210
rect 23378 30158 23390 30210
rect 27906 30158 27918 30210
rect 27970 30158 27982 30210
rect 20526 30146 20578 30158
rect 22766 30146 22818 30158
rect 27470 30146 27522 30158
rect 29150 30146 29202 30158
rect 29262 30210 29314 30222
rect 29262 30146 29314 30158
rect 30942 30210 30994 30222
rect 30942 30146 30994 30158
rect 31278 30210 31330 30222
rect 31278 30146 31330 30158
rect 33518 30210 33570 30222
rect 35634 30158 35646 30210
rect 35698 30158 35710 30210
rect 33518 30146 33570 30158
rect 6302 30098 6354 30110
rect 6302 30034 6354 30046
rect 6526 30098 6578 30110
rect 6526 30034 6578 30046
rect 7310 30098 7362 30110
rect 10558 30098 10610 30110
rect 9426 30046 9438 30098
rect 9490 30046 9502 30098
rect 7310 30034 7362 30046
rect 10558 30034 10610 30046
rect 12014 30098 12066 30110
rect 12014 30034 12066 30046
rect 12574 30098 12626 30110
rect 12574 30034 12626 30046
rect 16158 30098 16210 30110
rect 16158 30034 16210 30046
rect 17614 30098 17666 30110
rect 17614 30034 17666 30046
rect 20414 30098 20466 30110
rect 25006 30098 25058 30110
rect 27358 30098 27410 30110
rect 24210 30046 24222 30098
rect 24274 30046 24286 30098
rect 26338 30046 26350 30098
rect 26402 30046 26414 30098
rect 26898 30046 26910 30098
rect 26962 30046 26974 30098
rect 20414 30034 20466 30046
rect 25006 30034 25058 30046
rect 27358 30034 27410 30046
rect 30606 30098 30658 30110
rect 34974 30098 35026 30110
rect 31938 30046 31950 30098
rect 32002 30046 32014 30098
rect 30606 30034 30658 30046
rect 34974 30034 35026 30046
rect 5182 29986 5234 29998
rect 5182 29922 5234 29934
rect 6638 29986 6690 29998
rect 6638 29922 6690 29934
rect 14926 29986 14978 29998
rect 14926 29922 14978 29934
rect 20190 29986 20242 29998
rect 20190 29922 20242 29934
rect 20302 29986 20354 29998
rect 20302 29922 20354 29934
rect 22094 29986 22146 29998
rect 22094 29922 22146 29934
rect 25454 29986 25506 29998
rect 25454 29922 25506 29934
rect 25790 29986 25842 29998
rect 25790 29922 25842 29934
rect 29822 29986 29874 29998
rect 29822 29922 29874 29934
rect 30382 29986 30434 29998
rect 30382 29922 30434 29934
rect 31054 29986 31106 29998
rect 33954 29934 33966 29986
rect 34018 29934 34030 29986
rect 31054 29922 31106 29934
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 5742 29650 5794 29662
rect 5742 29586 5794 29598
rect 7086 29650 7138 29662
rect 7086 29586 7138 29598
rect 9102 29650 9154 29662
rect 9102 29586 9154 29598
rect 10222 29650 10274 29662
rect 10222 29586 10274 29598
rect 10446 29650 10498 29662
rect 10446 29586 10498 29598
rect 10894 29650 10946 29662
rect 17614 29650 17666 29662
rect 14578 29598 14590 29650
rect 14642 29598 14654 29650
rect 10894 29586 10946 29598
rect 17614 29586 17666 29598
rect 19406 29650 19458 29662
rect 19406 29586 19458 29598
rect 20414 29650 20466 29662
rect 20414 29586 20466 29598
rect 32062 29650 32114 29662
rect 32062 29586 32114 29598
rect 32510 29650 32562 29662
rect 32510 29586 32562 29598
rect 34526 29650 34578 29662
rect 34526 29586 34578 29598
rect 2046 29538 2098 29550
rect 2046 29474 2098 29486
rect 8430 29538 8482 29550
rect 8430 29474 8482 29486
rect 8766 29538 8818 29550
rect 8766 29474 8818 29486
rect 8878 29538 8930 29550
rect 8878 29474 8930 29486
rect 9886 29538 9938 29550
rect 15486 29538 15538 29550
rect 13682 29486 13694 29538
rect 13746 29486 13758 29538
rect 9886 29474 9938 29486
rect 15486 29474 15538 29486
rect 17502 29538 17554 29550
rect 17502 29474 17554 29486
rect 19070 29538 19122 29550
rect 19070 29474 19122 29486
rect 24334 29538 24386 29550
rect 24334 29474 24386 29486
rect 24670 29538 24722 29550
rect 31378 29486 31390 29538
rect 31442 29486 31454 29538
rect 24670 29474 24722 29486
rect 1710 29426 1762 29438
rect 1710 29362 1762 29374
rect 5630 29426 5682 29438
rect 5630 29362 5682 29374
rect 5854 29426 5906 29438
rect 7534 29426 7586 29438
rect 9774 29426 9826 29438
rect 6178 29374 6190 29426
rect 6242 29374 6254 29426
rect 7970 29374 7982 29426
rect 8034 29374 8046 29426
rect 5854 29362 5906 29374
rect 7534 29362 7586 29374
rect 9774 29362 9826 29374
rect 10110 29426 10162 29438
rect 10110 29362 10162 29374
rect 10558 29426 10610 29438
rect 16382 29426 16434 29438
rect 13570 29374 13582 29426
rect 13634 29374 13646 29426
rect 14690 29374 14702 29426
rect 14754 29374 14766 29426
rect 16146 29374 16158 29426
rect 16210 29374 16222 29426
rect 10558 29362 10610 29374
rect 16382 29362 16434 29374
rect 18174 29426 18226 29438
rect 19518 29426 19570 29438
rect 18610 29374 18622 29426
rect 18674 29374 18686 29426
rect 18174 29362 18226 29374
rect 19518 29362 19570 29374
rect 19630 29426 19682 29438
rect 19630 29362 19682 29374
rect 20078 29426 20130 29438
rect 20078 29362 20130 29374
rect 20302 29426 20354 29438
rect 33966 29426 34018 29438
rect 26338 29374 26350 29426
rect 26402 29374 26414 29426
rect 33506 29374 33518 29426
rect 33570 29374 33582 29426
rect 20302 29362 20354 29374
rect 33966 29362 34018 29374
rect 34750 29426 34802 29438
rect 34750 29362 34802 29374
rect 35198 29426 35250 29438
rect 35198 29362 35250 29374
rect 35422 29426 35474 29438
rect 38994 29374 39006 29426
rect 39058 29374 39070 29426
rect 35422 29362 35474 29374
rect 2494 29314 2546 29326
rect 2494 29250 2546 29262
rect 5294 29314 5346 29326
rect 6638 29314 6690 29326
rect 6178 29262 6190 29314
rect 6242 29311 6254 29314
rect 6402 29311 6414 29314
rect 6242 29265 6414 29311
rect 6242 29262 6254 29265
rect 6402 29262 6414 29265
rect 6466 29262 6478 29314
rect 5294 29250 5346 29262
rect 6638 29250 6690 29262
rect 11006 29314 11058 29326
rect 11006 29250 11058 29262
rect 20974 29314 21026 29326
rect 20974 29250 21026 29262
rect 25230 29314 25282 29326
rect 25230 29250 25282 29262
rect 25790 29314 25842 29326
rect 25790 29250 25842 29262
rect 33070 29314 33122 29326
rect 34974 29314 35026 29326
rect 34626 29262 34638 29314
rect 34690 29262 34702 29314
rect 33070 29250 33122 29262
rect 34974 29250 35026 29262
rect 35870 29314 35922 29326
rect 40114 29262 40126 29314
rect 40178 29262 40190 29314
rect 35870 29250 35922 29262
rect 17614 29202 17666 29214
rect 17614 29138 17666 29150
rect 20414 29202 20466 29214
rect 20414 29138 20466 29150
rect 25342 29202 25394 29214
rect 25342 29138 25394 29150
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 16718 28866 16770 28878
rect 11778 28814 11790 28866
rect 11842 28863 11854 28866
rect 12898 28863 12910 28866
rect 11842 28817 12910 28863
rect 11842 28814 11854 28817
rect 12898 28814 12910 28817
rect 12962 28814 12974 28866
rect 16718 28802 16770 28814
rect 17838 28866 17890 28878
rect 17838 28802 17890 28814
rect 26686 28866 26738 28878
rect 26686 28802 26738 28814
rect 31054 28866 31106 28878
rect 31054 28802 31106 28814
rect 32510 28866 32562 28878
rect 32510 28802 32562 28814
rect 8318 28754 8370 28766
rect 11902 28754 11954 28766
rect 9202 28702 9214 28754
rect 9266 28702 9278 28754
rect 10098 28702 10110 28754
rect 10162 28702 10174 28754
rect 8318 28690 8370 28702
rect 11902 28690 11954 28702
rect 12910 28754 12962 28766
rect 15486 28754 15538 28766
rect 14130 28702 14142 28754
rect 14194 28702 14206 28754
rect 12910 28690 12962 28702
rect 15486 28690 15538 28702
rect 16942 28754 16994 28766
rect 16942 28690 16994 28702
rect 17950 28754 18002 28766
rect 17950 28690 18002 28702
rect 19966 28754 20018 28766
rect 19966 28690 20018 28702
rect 21422 28754 21474 28766
rect 21422 28690 21474 28702
rect 21758 28754 21810 28766
rect 21758 28690 21810 28702
rect 27358 28754 27410 28766
rect 27358 28690 27410 28702
rect 27582 28754 27634 28766
rect 27582 28690 27634 28702
rect 27918 28754 27970 28766
rect 27918 28690 27970 28702
rect 28590 28754 28642 28766
rect 31502 28754 31554 28766
rect 29586 28702 29598 28754
rect 29650 28702 29662 28754
rect 28590 28690 28642 28702
rect 31502 28690 31554 28702
rect 33966 28754 34018 28766
rect 35522 28702 35534 28754
rect 35586 28702 35598 28754
rect 33966 28690 34018 28702
rect 2942 28642 2994 28654
rect 6638 28642 6690 28654
rect 6402 28590 6414 28642
rect 6466 28590 6478 28642
rect 2942 28578 2994 28590
rect 6638 28578 6690 28590
rect 6974 28642 7026 28654
rect 8206 28642 8258 28654
rect 11454 28642 11506 28654
rect 7634 28590 7646 28642
rect 7698 28590 7710 28642
rect 8978 28590 8990 28642
rect 9042 28590 9054 28642
rect 10434 28590 10446 28642
rect 10498 28590 10510 28642
rect 6974 28578 7026 28590
rect 8206 28578 8258 28590
rect 11454 28578 11506 28590
rect 12462 28642 12514 28654
rect 15150 28642 15202 28654
rect 17390 28642 17442 28654
rect 13570 28590 13582 28642
rect 13634 28590 13646 28642
rect 15922 28590 15934 28642
rect 15986 28590 15998 28642
rect 12462 28578 12514 28590
rect 15150 28578 15202 28590
rect 17390 28578 17442 28590
rect 22654 28642 22706 28654
rect 22654 28578 22706 28590
rect 22990 28642 23042 28654
rect 29150 28642 29202 28654
rect 23650 28590 23662 28642
rect 23714 28590 23726 28642
rect 22990 28578 23042 28590
rect 29150 28578 29202 28590
rect 30382 28642 30434 28654
rect 30382 28578 30434 28590
rect 31278 28642 31330 28654
rect 31278 28578 31330 28590
rect 31726 28642 31778 28654
rect 31726 28578 31778 28590
rect 31950 28642 32002 28654
rect 34302 28642 34354 28654
rect 33506 28590 33518 28642
rect 33570 28590 33582 28642
rect 31950 28578 32002 28590
rect 34302 28578 34354 28590
rect 34750 28642 34802 28654
rect 37102 28642 37154 28654
rect 35410 28590 35422 28642
rect 35474 28590 35486 28642
rect 36306 28590 36318 28642
rect 36370 28590 36382 28642
rect 34750 28578 34802 28590
rect 37102 28578 37154 28590
rect 37550 28642 37602 28654
rect 37550 28578 37602 28590
rect 39678 28642 39730 28654
rect 39678 28578 39730 28590
rect 40238 28642 40290 28654
rect 40238 28578 40290 28590
rect 6862 28530 6914 28542
rect 6862 28466 6914 28478
rect 9662 28530 9714 28542
rect 9662 28466 9714 28478
rect 11006 28530 11058 28542
rect 17278 28530 17330 28542
rect 13682 28478 13694 28530
rect 13746 28478 13758 28530
rect 16258 28478 16270 28530
rect 16322 28478 16334 28530
rect 11006 28466 11058 28478
rect 17278 28466 17330 28478
rect 25902 28530 25954 28542
rect 25902 28466 25954 28478
rect 27022 28530 27074 28542
rect 27022 28466 27074 28478
rect 27806 28530 27858 28542
rect 27806 28466 27858 28478
rect 28030 28530 28082 28542
rect 28030 28466 28082 28478
rect 32398 28530 32450 28542
rect 32398 28466 32450 28478
rect 32510 28530 32562 28542
rect 39902 28530 39954 28542
rect 33394 28478 33406 28530
rect 33458 28478 33470 28530
rect 32510 28466 32562 28478
rect 39902 28466 39954 28478
rect 2158 28418 2210 28430
rect 2158 28354 2210 28366
rect 5854 28418 5906 28430
rect 5854 28354 5906 28366
rect 5966 28418 6018 28430
rect 5966 28354 6018 28366
rect 6078 28418 6130 28430
rect 6078 28354 6130 28366
rect 17166 28418 17218 28430
rect 17166 28354 17218 28366
rect 18398 28418 18450 28430
rect 18398 28354 18450 28366
rect 19070 28418 19122 28430
rect 19070 28354 19122 28366
rect 21870 28418 21922 28430
rect 21870 28354 21922 28366
rect 31838 28418 31890 28430
rect 31838 28354 31890 28366
rect 36094 28418 36146 28430
rect 36094 28354 36146 28366
rect 36990 28418 37042 28430
rect 36990 28354 37042 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 7310 28082 7362 28094
rect 6738 28030 6750 28082
rect 6802 28030 6814 28082
rect 7310 28018 7362 28030
rect 7534 28082 7586 28094
rect 7534 28018 7586 28030
rect 8766 28082 8818 28094
rect 8766 28018 8818 28030
rect 10334 28082 10386 28094
rect 10334 28018 10386 28030
rect 10446 28082 10498 28094
rect 10446 28018 10498 28030
rect 10558 28082 10610 28094
rect 16606 28082 16658 28094
rect 14690 28030 14702 28082
rect 14754 28030 14766 28082
rect 10558 28018 10610 28030
rect 16606 28018 16658 28030
rect 17726 28082 17778 28094
rect 22542 28082 22594 28094
rect 21746 28030 21758 28082
rect 21810 28030 21822 28082
rect 17726 28018 17778 28030
rect 22542 28018 22594 28030
rect 22766 28082 22818 28094
rect 22766 28018 22818 28030
rect 23774 28082 23826 28094
rect 23774 28018 23826 28030
rect 24334 28082 24386 28094
rect 24334 28018 24386 28030
rect 26350 28082 26402 28094
rect 30718 28082 30770 28094
rect 29698 28030 29710 28082
rect 29762 28030 29774 28082
rect 26350 28018 26402 28030
rect 30718 28018 30770 28030
rect 32958 28082 33010 28094
rect 32958 28018 33010 28030
rect 33182 28082 33234 28094
rect 37438 28082 37490 28094
rect 36866 28030 36878 28082
rect 36930 28030 36942 28082
rect 33182 28018 33234 28030
rect 37438 28018 37490 28030
rect 8654 27970 8706 27982
rect 8654 27906 8706 27918
rect 23550 27970 23602 27982
rect 23550 27906 23602 27918
rect 23886 27970 23938 27982
rect 23886 27906 23938 27918
rect 30830 27970 30882 27982
rect 30830 27906 30882 27918
rect 33294 27970 33346 27982
rect 33294 27906 33346 27918
rect 3838 27858 3890 27870
rect 10222 27858 10274 27870
rect 19070 27858 19122 27870
rect 22990 27858 23042 27870
rect 4274 27806 4286 27858
rect 4338 27806 4350 27858
rect 10770 27806 10782 27858
rect 10834 27806 10846 27858
rect 11778 27806 11790 27858
rect 11842 27806 11854 27858
rect 12226 27806 12238 27858
rect 12290 27806 12302 27858
rect 19506 27806 19518 27858
rect 19570 27806 19582 27858
rect 3838 27794 3890 27806
rect 10222 27794 10274 27806
rect 19070 27794 19122 27806
rect 22990 27794 23042 27806
rect 23438 27858 23490 27870
rect 23438 27794 23490 27806
rect 26574 27858 26626 27870
rect 30382 27858 30434 27870
rect 33742 27858 33794 27870
rect 27234 27806 27246 27858
rect 27298 27806 27310 27858
rect 31938 27806 31950 27858
rect 32002 27806 32014 27858
rect 34402 27806 34414 27858
rect 34466 27806 34478 27858
rect 26574 27794 26626 27806
rect 30382 27794 30434 27806
rect 33742 27794 33794 27806
rect 7646 27746 7698 27758
rect 7646 27682 7698 27694
rect 8094 27746 8146 27758
rect 8094 27682 8146 27694
rect 11454 27746 11506 27758
rect 11454 27682 11506 27694
rect 15934 27746 15986 27758
rect 15934 27682 15986 27694
rect 22878 27746 22930 27758
rect 22878 27682 22930 27694
rect 25342 27746 25394 27758
rect 25342 27682 25394 27694
rect 31502 27746 31554 27758
rect 32274 27694 32286 27746
rect 32338 27694 32350 27746
rect 31502 27682 31554 27694
rect 15374 27634 15426 27646
rect 15374 27570 15426 27582
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 10446 27298 10498 27310
rect 10446 27234 10498 27246
rect 17054 27298 17106 27310
rect 17054 27234 17106 27246
rect 29598 27298 29650 27310
rect 30706 27246 30718 27298
rect 30770 27295 30782 27298
rect 31490 27295 31502 27298
rect 30770 27249 31502 27295
rect 30770 27246 30782 27249
rect 31490 27246 31502 27249
rect 31554 27246 31566 27298
rect 31714 27246 31726 27298
rect 31778 27246 31790 27298
rect 33842 27246 33854 27298
rect 33906 27295 33918 27298
rect 35186 27295 35198 27298
rect 33906 27249 35198 27295
rect 33906 27246 33918 27249
rect 35186 27246 35198 27249
rect 35250 27246 35262 27298
rect 29598 27234 29650 27246
rect 7422 27186 7474 27198
rect 12238 27186 12290 27198
rect 10770 27134 10782 27186
rect 10834 27134 10846 27186
rect 7422 27122 7474 27134
rect 12238 27122 12290 27134
rect 25454 27186 25506 27198
rect 27470 27186 27522 27198
rect 26674 27134 26686 27186
rect 26738 27134 26750 27186
rect 25454 27122 25506 27134
rect 27470 27122 27522 27134
rect 28590 27186 28642 27198
rect 28590 27122 28642 27134
rect 33406 27186 33458 27198
rect 33406 27122 33458 27134
rect 33854 27186 33906 27198
rect 33854 27122 33906 27134
rect 34750 27186 34802 27198
rect 34750 27122 34802 27134
rect 35198 27186 35250 27198
rect 35198 27122 35250 27134
rect 13358 27074 13410 27086
rect 19406 27074 19458 27086
rect 14018 27022 14030 27074
rect 14082 27022 14094 27074
rect 18274 27022 18286 27074
rect 18338 27022 18350 27074
rect 13358 27010 13410 27022
rect 19406 27010 19458 27022
rect 21198 27074 21250 27086
rect 25006 27074 25058 27086
rect 21858 27022 21870 27074
rect 21922 27022 21934 27074
rect 21198 27010 21250 27022
rect 25006 27010 25058 27022
rect 25902 27074 25954 27086
rect 25902 27010 25954 27022
rect 26238 27074 26290 27086
rect 26238 27010 26290 27022
rect 30942 27074 30994 27086
rect 30942 27010 30994 27022
rect 32174 27074 32226 27086
rect 32498 27022 32510 27074
rect 32562 27022 32574 27074
rect 32174 27010 32226 27022
rect 8430 26962 8482 26974
rect 8430 26898 8482 26910
rect 10670 26962 10722 26974
rect 10670 26898 10722 26910
rect 11118 26962 11170 26974
rect 11118 26898 11170 26910
rect 11230 26962 11282 26974
rect 11230 26898 11282 26910
rect 12350 26962 12402 26974
rect 27806 26962 27858 26974
rect 17378 26910 17390 26962
rect 17442 26910 17454 26962
rect 12350 26898 12402 26910
rect 27806 26898 27858 26910
rect 28142 26962 28194 26974
rect 28142 26898 28194 26910
rect 29262 26962 29314 26974
rect 32286 26962 32338 26974
rect 29810 26910 29822 26962
rect 29874 26910 29886 26962
rect 30370 26910 30382 26962
rect 30434 26910 30446 26962
rect 29262 26898 29314 26910
rect 32286 26898 32338 26910
rect 10222 26850 10274 26862
rect 10222 26786 10274 26798
rect 11342 26850 11394 26862
rect 11342 26786 11394 26798
rect 12126 26850 12178 26862
rect 12126 26786 12178 26798
rect 12574 26850 12626 26862
rect 18958 26850 19010 26862
rect 31390 26850 31442 26862
rect 16258 26798 16270 26850
rect 16322 26798 16334 26850
rect 24098 26798 24110 26850
rect 24162 26798 24174 26850
rect 12574 26786 12626 26798
rect 18958 26786 19010 26798
rect 31390 26786 31442 26798
rect 33070 26850 33122 26862
rect 33070 26786 33122 26798
rect 34302 26850 34354 26862
rect 34302 26786 34354 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 6414 26514 6466 26526
rect 6414 26450 6466 26462
rect 7758 26514 7810 26526
rect 7758 26450 7810 26462
rect 16046 26514 16098 26526
rect 16046 26450 16098 26462
rect 23102 26514 23154 26526
rect 23102 26450 23154 26462
rect 23886 26514 23938 26526
rect 34414 26514 34466 26526
rect 33394 26462 33406 26514
rect 33458 26462 33470 26514
rect 23886 26450 23938 26462
rect 34414 26450 34466 26462
rect 7534 26402 7586 26414
rect 7534 26338 7586 26350
rect 8654 26402 8706 26414
rect 23214 26402 23266 26414
rect 13346 26350 13358 26402
rect 13410 26350 13422 26402
rect 8654 26338 8706 26350
rect 23214 26338 23266 26350
rect 31950 26402 32002 26414
rect 31950 26338 32002 26350
rect 32510 26402 32562 26414
rect 32510 26338 32562 26350
rect 7982 26290 8034 26302
rect 2818 26238 2830 26290
rect 2882 26238 2894 26290
rect 7982 26226 8034 26238
rect 8094 26290 8146 26302
rect 8094 26226 8146 26238
rect 8542 26290 8594 26302
rect 8542 26226 8594 26238
rect 8878 26290 8930 26302
rect 8878 26226 8930 26238
rect 9662 26290 9714 26302
rect 15934 26290 15986 26302
rect 15474 26238 15486 26290
rect 15538 26238 15550 26290
rect 9662 26226 9714 26238
rect 15934 26226 15986 26238
rect 16494 26290 16546 26302
rect 19966 26290 20018 26302
rect 22430 26290 22482 26302
rect 22990 26290 23042 26302
rect 26350 26290 26402 26302
rect 29038 26290 29090 26302
rect 18498 26238 18510 26290
rect 18562 26238 18574 26290
rect 21970 26238 21982 26290
rect 22034 26238 22046 26290
rect 22754 26238 22766 26290
rect 22818 26238 22830 26290
rect 23426 26238 23438 26290
rect 23490 26238 23502 26290
rect 26674 26238 26686 26290
rect 26738 26238 26750 26290
rect 16494 26226 16546 26238
rect 19966 26226 20018 26238
rect 22430 26226 22482 26238
rect 22990 26226 23042 26238
rect 26350 26226 26402 26238
rect 29038 26226 29090 26238
rect 29486 26290 29538 26302
rect 29486 26226 29538 26238
rect 29710 26290 29762 26302
rect 29710 26226 29762 26238
rect 31166 26290 31218 26302
rect 31166 26226 31218 26238
rect 32174 26290 32226 26302
rect 32174 26226 32226 26238
rect 32958 26290 33010 26302
rect 33966 26290 34018 26302
rect 33282 26238 33294 26290
rect 33346 26238 33358 26290
rect 38994 26238 39006 26290
rect 39058 26238 39070 26290
rect 32958 26226 33010 26238
rect 33966 26226 34018 26238
rect 6974 26178 7026 26190
rect 1922 26126 1934 26178
rect 1986 26126 1998 26178
rect 6974 26114 7026 26126
rect 7870 26178 7922 26190
rect 19294 26178 19346 26190
rect 23774 26178 23826 26190
rect 17938 26126 17950 26178
rect 18002 26126 18014 26178
rect 18610 26126 18622 26178
rect 18674 26175 18686 26178
rect 19058 26175 19070 26178
rect 18674 26129 19070 26175
rect 18674 26126 18686 26129
rect 19058 26126 19070 26129
rect 19122 26126 19134 26178
rect 21522 26126 21534 26178
rect 21586 26126 21598 26178
rect 7870 26114 7922 26126
rect 19294 26114 19346 26126
rect 23774 26114 23826 26126
rect 24334 26178 24386 26190
rect 28478 26178 28530 26190
rect 27346 26126 27358 26178
rect 27410 26126 27422 26178
rect 24334 26114 24386 26126
rect 28478 26114 28530 26126
rect 28814 26178 28866 26190
rect 28814 26114 28866 26126
rect 29262 26178 29314 26190
rect 30718 26178 30770 26190
rect 30370 26126 30382 26178
rect 30434 26126 30446 26178
rect 29262 26114 29314 26126
rect 30718 26114 30770 26126
rect 31614 26178 31666 26190
rect 31614 26114 31666 26126
rect 32062 26178 32114 26190
rect 32062 26114 32114 26126
rect 33742 26178 33794 26190
rect 33742 26114 33794 26126
rect 34862 26178 34914 26190
rect 34862 26114 34914 26126
rect 35310 26178 35362 26190
rect 40114 26126 40126 26178
rect 40178 26126 40190 26178
rect 35310 26114 35362 26126
rect 19406 26066 19458 26078
rect 19406 26002 19458 26014
rect 33518 26066 33570 26078
rect 33518 26002 33570 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 8766 25730 8818 25742
rect 8766 25666 8818 25678
rect 13582 25730 13634 25742
rect 13582 25666 13634 25678
rect 14702 25730 14754 25742
rect 14702 25666 14754 25678
rect 20302 25730 20354 25742
rect 20302 25666 20354 25678
rect 21534 25730 21586 25742
rect 21534 25666 21586 25678
rect 36542 25730 36594 25742
rect 36542 25666 36594 25678
rect 7310 25618 7362 25630
rect 12574 25618 12626 25630
rect 10434 25566 10446 25618
rect 10498 25566 10510 25618
rect 12114 25566 12126 25618
rect 12178 25566 12190 25618
rect 7310 25554 7362 25566
rect 12574 25554 12626 25566
rect 12686 25618 12738 25630
rect 12686 25554 12738 25566
rect 14814 25618 14866 25630
rect 14814 25554 14866 25566
rect 15262 25618 15314 25630
rect 15262 25554 15314 25566
rect 16382 25618 16434 25630
rect 16382 25554 16434 25566
rect 23774 25618 23826 25630
rect 23774 25554 23826 25566
rect 24222 25618 24274 25630
rect 24222 25554 24274 25566
rect 2942 25506 2994 25518
rect 2942 25442 2994 25454
rect 4734 25506 4786 25518
rect 4734 25442 4786 25454
rect 5070 25506 5122 25518
rect 5070 25442 5122 25454
rect 5630 25506 5682 25518
rect 5630 25442 5682 25454
rect 5854 25506 5906 25518
rect 6414 25506 6466 25518
rect 6178 25454 6190 25506
rect 6242 25454 6254 25506
rect 5854 25442 5906 25454
rect 6414 25442 6466 25454
rect 6750 25506 6802 25518
rect 8206 25506 8258 25518
rect 7970 25454 7982 25506
rect 8034 25454 8046 25506
rect 6750 25442 6802 25454
rect 8206 25442 8258 25454
rect 9438 25506 9490 25518
rect 9438 25442 9490 25454
rect 9774 25506 9826 25518
rect 12014 25506 12066 25518
rect 10322 25454 10334 25506
rect 10386 25454 10398 25506
rect 11554 25454 11566 25506
rect 11618 25454 11630 25506
rect 9774 25442 9826 25454
rect 12014 25442 12066 25454
rect 13694 25506 13746 25518
rect 13694 25442 13746 25454
rect 14366 25506 14418 25518
rect 14366 25442 14418 25454
rect 16606 25506 16658 25518
rect 22430 25506 22482 25518
rect 24782 25506 24834 25518
rect 29822 25506 29874 25518
rect 31502 25506 31554 25518
rect 17266 25454 17278 25506
rect 17330 25454 17342 25506
rect 22866 25454 22878 25506
rect 22930 25454 22942 25506
rect 25218 25454 25230 25506
rect 25282 25454 25294 25506
rect 29586 25454 29598 25506
rect 29650 25454 29662 25506
rect 30034 25454 30046 25506
rect 30098 25454 30110 25506
rect 30818 25454 30830 25506
rect 30882 25454 30894 25506
rect 16606 25442 16658 25454
rect 22430 25442 22482 25454
rect 24782 25442 24834 25454
rect 29822 25442 29874 25454
rect 31502 25442 31554 25454
rect 32846 25506 32898 25518
rect 39006 25506 39058 25518
rect 33394 25454 33406 25506
rect 33458 25454 33470 25506
rect 32846 25442 32898 25454
rect 39006 25442 39058 25454
rect 8654 25394 8706 25406
rect 8654 25330 8706 25342
rect 9550 25394 9602 25406
rect 9550 25330 9602 25342
rect 11230 25394 11282 25406
rect 11230 25330 11282 25342
rect 12126 25394 12178 25406
rect 12126 25330 12178 25342
rect 13582 25394 13634 25406
rect 13582 25330 13634 25342
rect 14030 25394 14082 25406
rect 14030 25330 14082 25342
rect 19518 25394 19570 25406
rect 19518 25330 19570 25342
rect 21422 25394 21474 25406
rect 21422 25330 21474 25342
rect 23326 25394 23378 25406
rect 23326 25330 23378 25342
rect 30270 25394 30322 25406
rect 30270 25330 30322 25342
rect 31726 25394 31778 25406
rect 31726 25330 31778 25342
rect 2158 25282 2210 25294
rect 2158 25218 2210 25230
rect 4958 25282 5010 25294
rect 4958 25218 5010 25230
rect 5742 25282 5794 25294
rect 5742 25218 5794 25230
rect 6638 25282 6690 25294
rect 6638 25218 6690 25230
rect 8766 25282 8818 25294
rect 8766 25218 8818 25230
rect 11790 25282 11842 25294
rect 11790 25218 11842 25230
rect 12798 25282 12850 25294
rect 12798 25218 12850 25230
rect 15710 25282 15762 25294
rect 15710 25218 15762 25230
rect 20638 25282 20690 25294
rect 20638 25218 20690 25230
rect 21534 25282 21586 25294
rect 28254 25282 28306 25294
rect 27458 25230 27470 25282
rect 27522 25230 27534 25282
rect 21534 25218 21586 25230
rect 28254 25218 28306 25230
rect 28590 25282 28642 25294
rect 32062 25282 32114 25294
rect 29810 25230 29822 25282
rect 29874 25230 29886 25282
rect 28590 25218 28642 25230
rect 32062 25218 32114 25230
rect 32174 25282 32226 25294
rect 32174 25218 32226 25230
rect 32286 25282 32338 25294
rect 32286 25218 32338 25230
rect 32510 25282 32562 25294
rect 39790 25282 39842 25294
rect 35970 25230 35982 25282
rect 36034 25230 36046 25282
rect 32510 25218 32562 25230
rect 39790 25218 39842 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 2830 24946 2882 24958
rect 6862 24946 6914 24958
rect 2034 24894 2046 24946
rect 2098 24894 2110 24946
rect 3602 24894 3614 24946
rect 3666 24894 3678 24946
rect 2830 24882 2882 24894
rect 6862 24882 6914 24894
rect 10110 24946 10162 24958
rect 10110 24882 10162 24894
rect 10222 24946 10274 24958
rect 10222 24882 10274 24894
rect 13806 24946 13858 24958
rect 13806 24882 13858 24894
rect 15822 24946 15874 24958
rect 15822 24882 15874 24894
rect 18734 24946 18786 24958
rect 18734 24882 18786 24894
rect 18846 24946 18898 24958
rect 18846 24882 18898 24894
rect 19630 24946 19682 24958
rect 19630 24882 19682 24894
rect 20302 24946 20354 24958
rect 20302 24882 20354 24894
rect 21198 24946 21250 24958
rect 21198 24882 21250 24894
rect 24446 24946 24498 24958
rect 24446 24882 24498 24894
rect 25454 24946 25506 24958
rect 25454 24882 25506 24894
rect 25902 24946 25954 24958
rect 25902 24882 25954 24894
rect 26686 24946 26738 24958
rect 26686 24882 26738 24894
rect 26798 24946 26850 24958
rect 26798 24882 26850 24894
rect 27358 24946 27410 24958
rect 27358 24882 27410 24894
rect 35982 24946 36034 24958
rect 35982 24882 36034 24894
rect 36654 24946 36706 24958
rect 36654 24882 36706 24894
rect 7982 24834 8034 24846
rect 7982 24770 8034 24782
rect 9550 24834 9602 24846
rect 9550 24770 9602 24782
rect 10446 24834 10498 24846
rect 17502 24834 17554 24846
rect 11330 24782 11342 24834
rect 11394 24782 11406 24834
rect 15250 24782 15262 24834
rect 15314 24782 15326 24834
rect 10446 24770 10498 24782
rect 17502 24770 17554 24782
rect 19406 24834 19458 24846
rect 19406 24770 19458 24782
rect 19742 24834 19794 24846
rect 19742 24770 19794 24782
rect 20526 24834 20578 24846
rect 20526 24770 20578 24782
rect 22654 24834 22706 24846
rect 22654 24770 22706 24782
rect 22990 24834 23042 24846
rect 22990 24770 23042 24782
rect 23774 24834 23826 24846
rect 23774 24770 23826 24782
rect 25790 24834 25842 24846
rect 25790 24770 25842 24782
rect 26126 24834 26178 24846
rect 26126 24770 26178 24782
rect 27246 24834 27298 24846
rect 27246 24770 27298 24782
rect 30494 24834 30546 24846
rect 30494 24770 30546 24782
rect 31502 24834 31554 24846
rect 31502 24770 31554 24782
rect 33070 24834 33122 24846
rect 33070 24770 33122 24782
rect 33182 24834 33234 24846
rect 33182 24770 33234 24782
rect 36206 24834 36258 24846
rect 36206 24770 36258 24782
rect 1710 24722 1762 24734
rect 6526 24722 6578 24734
rect 9998 24722 10050 24734
rect 17390 24722 17442 24734
rect 5842 24670 5854 24722
rect 5906 24670 5918 24722
rect 8418 24670 8430 24722
rect 8482 24670 8494 24722
rect 11218 24670 11230 24722
rect 11282 24670 11294 24722
rect 12898 24670 12910 24722
rect 12962 24670 12974 24722
rect 14914 24670 14926 24722
rect 14978 24670 14990 24722
rect 1710 24658 1762 24670
rect 6526 24658 6578 24670
rect 9998 24658 10050 24670
rect 17390 24658 17442 24670
rect 17726 24722 17778 24734
rect 17726 24658 17778 24670
rect 18622 24722 18674 24734
rect 18622 24658 18674 24670
rect 19294 24722 19346 24734
rect 19294 24658 19346 24670
rect 20190 24722 20242 24734
rect 21086 24722 21138 24734
rect 20738 24670 20750 24722
rect 20802 24670 20814 24722
rect 20190 24658 20242 24670
rect 21086 24658 21138 24670
rect 21310 24722 21362 24734
rect 23998 24722 24050 24734
rect 22082 24670 22094 24722
rect 22146 24670 22158 24722
rect 23314 24670 23326 24722
rect 23378 24670 23390 24722
rect 21310 24658 21362 24670
rect 23998 24658 24050 24670
rect 24334 24722 24386 24734
rect 24334 24658 24386 24670
rect 26238 24722 26290 24734
rect 26238 24658 26290 24670
rect 26910 24722 26962 24734
rect 26910 24658 26962 24670
rect 27582 24722 27634 24734
rect 36318 24722 36370 24734
rect 28242 24670 28254 24722
rect 28306 24670 28318 24722
rect 31714 24670 31726 24722
rect 31778 24670 31790 24722
rect 32162 24670 32174 24722
rect 32226 24670 32238 24722
rect 34290 24670 34302 24722
rect 34354 24670 34366 24722
rect 35634 24670 35646 24722
rect 35698 24670 35710 24722
rect 27582 24658 27634 24670
rect 36318 24658 36370 24670
rect 2494 24610 2546 24622
rect 16382 24610 16434 24622
rect 8866 24558 8878 24610
rect 8930 24558 8942 24610
rect 2494 24546 2546 24558
rect 16382 24546 16434 24558
rect 16830 24610 16882 24622
rect 16830 24546 16882 24558
rect 18062 24610 18114 24622
rect 31278 24610 31330 24622
rect 36766 24610 36818 24622
rect 22194 24558 22206 24610
rect 22258 24558 22270 24610
rect 23202 24558 23214 24610
rect 23266 24558 23278 24610
rect 23650 24558 23662 24610
rect 23714 24558 23726 24610
rect 34402 24558 34414 24610
rect 34466 24558 34478 24610
rect 35410 24558 35422 24610
rect 35474 24558 35486 24610
rect 18062 24546 18114 24558
rect 31278 24546 31330 24558
rect 36766 24546 36818 24558
rect 37214 24610 37266 24622
rect 37214 24546 37266 24558
rect 9662 24498 9714 24510
rect 9662 24434 9714 24446
rect 17950 24498 18002 24510
rect 17950 24434 18002 24446
rect 24446 24498 24498 24510
rect 24446 24434 24498 24446
rect 33182 24498 33234 24510
rect 34178 24446 34190 24498
rect 34242 24446 34254 24498
rect 33182 24434 33234 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 9214 24162 9266 24174
rect 29598 24162 29650 24174
rect 28466 24110 28478 24162
rect 28530 24110 28542 24162
rect 9214 24098 9266 24110
rect 29598 24098 29650 24110
rect 8542 24050 8594 24062
rect 10670 24050 10722 24062
rect 14478 24050 14530 24062
rect 7634 23998 7646 24050
rect 7698 23998 7710 24050
rect 9538 23998 9550 24050
rect 9602 23998 9614 24050
rect 13682 23998 13694 24050
rect 13746 23998 13758 24050
rect 8542 23986 8594 23998
rect 10670 23986 10722 23998
rect 14478 23986 14530 23998
rect 19406 24050 19458 24062
rect 27134 24050 27186 24062
rect 20290 23998 20302 24050
rect 20354 23998 20366 24050
rect 21746 23998 21758 24050
rect 21810 23998 21822 24050
rect 19406 23986 19458 23998
rect 27134 23986 27186 23998
rect 29486 24050 29538 24062
rect 29486 23986 29538 23998
rect 33966 24050 34018 24062
rect 40002 23998 40014 24050
rect 40066 23998 40078 24050
rect 33966 23986 34018 23998
rect 2270 23938 2322 23950
rect 2270 23874 2322 23886
rect 7086 23938 7138 23950
rect 7086 23874 7138 23886
rect 7198 23938 7250 23950
rect 10334 23938 10386 23950
rect 14702 23938 14754 23950
rect 25006 23938 25058 23950
rect 28254 23938 28306 23950
rect 8082 23886 8094 23938
rect 8146 23886 8158 23938
rect 10546 23886 10558 23938
rect 10610 23886 10622 23938
rect 12002 23886 12014 23938
rect 12066 23886 12078 23938
rect 12562 23886 12574 23938
rect 12626 23886 12638 23938
rect 15362 23886 15374 23938
rect 15426 23886 15438 23938
rect 20066 23886 20078 23938
rect 20130 23886 20142 23938
rect 22418 23886 22430 23938
rect 22482 23886 22494 23938
rect 23986 23886 23998 23938
rect 24050 23886 24062 23938
rect 25890 23886 25902 23938
rect 25954 23886 25966 23938
rect 7198 23874 7250 23886
rect 10334 23874 10386 23886
rect 14702 23874 14754 23886
rect 25006 23874 25058 23886
rect 28254 23874 28306 23886
rect 28366 23938 28418 23950
rect 35422 23938 35474 23950
rect 30370 23886 30382 23938
rect 30434 23886 30446 23938
rect 33058 23886 33070 23938
rect 33122 23886 33134 23938
rect 33506 23886 33518 23938
rect 33570 23886 33582 23938
rect 34178 23886 34190 23938
rect 34242 23886 34254 23938
rect 34626 23886 34638 23938
rect 34690 23886 34702 23938
rect 28366 23874 28418 23886
rect 35422 23874 35474 23886
rect 35870 23938 35922 23950
rect 38994 23886 39006 23938
rect 39058 23886 39070 23938
rect 35870 23874 35922 23886
rect 9438 23826 9490 23838
rect 13470 23826 13522 23838
rect 11106 23774 11118 23826
rect 11170 23774 11182 23826
rect 9438 23762 9490 23774
rect 13470 23762 13522 23774
rect 18734 23826 18786 23838
rect 18734 23762 18786 23774
rect 20750 23826 20802 23838
rect 20750 23762 20802 23774
rect 21310 23826 21362 23838
rect 26798 23826 26850 23838
rect 22978 23774 22990 23826
rect 23042 23774 23054 23826
rect 30482 23774 30494 23826
rect 30546 23774 30558 23826
rect 21310 23762 21362 23774
rect 26798 23762 26850 23774
rect 1710 23714 1762 23726
rect 1710 23650 1762 23662
rect 2718 23714 2770 23726
rect 18398 23714 18450 23726
rect 17826 23662 17838 23714
rect 17890 23662 17902 23714
rect 2718 23650 2770 23662
rect 18398 23650 18450 23662
rect 21534 23714 21586 23726
rect 21534 23650 21586 23662
rect 21758 23714 21810 23726
rect 21758 23650 21810 23662
rect 21870 23714 21922 23726
rect 27022 23714 27074 23726
rect 23314 23662 23326 23714
rect 23378 23662 23390 23714
rect 21870 23650 21922 23662
rect 27022 23650 27074 23662
rect 27246 23714 27298 23726
rect 27246 23650 27298 23662
rect 27358 23714 27410 23726
rect 31154 23662 31166 23714
rect 31218 23662 31230 23714
rect 27358 23650 27410 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 3390 23378 3442 23390
rect 3390 23314 3442 23326
rect 5406 23378 5458 23390
rect 5406 23314 5458 23326
rect 16270 23378 16322 23390
rect 16270 23314 16322 23326
rect 18398 23378 18450 23390
rect 18398 23314 18450 23326
rect 19630 23378 19682 23390
rect 19630 23314 19682 23326
rect 20078 23378 20130 23390
rect 21198 23378 21250 23390
rect 34862 23378 34914 23390
rect 20962 23326 20974 23378
rect 21026 23326 21038 23378
rect 22978 23326 22990 23378
rect 23042 23326 23054 23378
rect 27346 23326 27358 23378
rect 27410 23326 27422 23378
rect 33282 23326 33294 23378
rect 33346 23326 33358 23378
rect 20078 23314 20130 23326
rect 21198 23314 21250 23326
rect 34862 23314 34914 23326
rect 39006 23378 39058 23390
rect 39006 23314 39058 23326
rect 8654 23266 8706 23278
rect 12126 23266 12178 23278
rect 7298 23214 7310 23266
rect 7362 23214 7374 23266
rect 9650 23214 9662 23266
rect 9714 23214 9726 23266
rect 8654 23202 8706 23214
rect 12126 23202 12178 23214
rect 17502 23266 17554 23278
rect 26686 23266 26738 23278
rect 34638 23266 34690 23278
rect 39902 23266 39954 23278
rect 25218 23214 25230 23266
rect 25282 23214 25294 23266
rect 34066 23214 34078 23266
rect 34130 23214 34142 23266
rect 39218 23214 39230 23266
rect 39282 23214 39294 23266
rect 17502 23202 17554 23214
rect 8318 23154 8370 23166
rect 2818 23102 2830 23154
rect 2882 23102 2894 23154
rect 8318 23090 8370 23102
rect 8766 23154 8818 23166
rect 16158 23154 16210 23166
rect 9538 23102 9550 23154
rect 9602 23102 9614 23154
rect 11554 23102 11566 23154
rect 11618 23102 11630 23154
rect 8766 23090 8818 23102
rect 16158 23090 16210 23102
rect 17390 23154 17442 23166
rect 17390 23090 17442 23102
rect 17614 23154 17666 23166
rect 20414 23154 20466 23166
rect 17938 23102 17950 23154
rect 18002 23102 18014 23154
rect 17614 23090 17666 23102
rect 20414 23090 20466 23102
rect 20638 23154 20690 23166
rect 22082 23158 22094 23210
rect 22146 23158 22158 23210
rect 26686 23202 26738 23214
rect 34638 23202 34690 23214
rect 39902 23202 39954 23214
rect 20638 23090 20690 23102
rect 22430 23154 22482 23166
rect 22430 23090 22482 23102
rect 22654 23154 22706 23166
rect 24558 23154 24610 23166
rect 26462 23154 26514 23166
rect 24210 23102 24222 23154
rect 24274 23102 24286 23154
rect 25442 23102 25454 23154
rect 25506 23102 25518 23154
rect 25890 23102 25902 23154
rect 25954 23102 25966 23154
rect 22654 23090 22706 23102
rect 24558 23090 24610 23102
rect 26462 23090 26514 23102
rect 26798 23154 26850 23166
rect 26798 23090 26850 23102
rect 27918 23154 27970 23166
rect 31390 23154 31442 23166
rect 34526 23154 34578 23166
rect 28578 23102 28590 23154
rect 28642 23102 28654 23154
rect 32162 23102 32174 23154
rect 32226 23102 32238 23154
rect 33170 23102 33182 23154
rect 33234 23102 33246 23154
rect 33954 23102 33966 23154
rect 34018 23102 34030 23154
rect 27918 23090 27970 23102
rect 31390 23090 31442 23102
rect 34526 23090 34578 23102
rect 39566 23154 39618 23166
rect 39566 23090 39618 23102
rect 40238 23154 40290 23166
rect 40238 23090 40290 23102
rect 8430 23042 8482 23054
rect 16830 23042 16882 23054
rect 1922 22990 1934 23042
rect 1986 22990 1998 23042
rect 11442 22990 11454 23042
rect 11506 22990 11518 23042
rect 8430 22978 8482 22990
rect 16830 22978 16882 22990
rect 19294 23042 19346 23054
rect 19294 22978 19346 22990
rect 19966 23042 20018 23054
rect 19966 22978 20018 22990
rect 21870 23042 21922 23054
rect 21870 22978 21922 22990
rect 24670 23042 24722 23054
rect 24670 22978 24722 22990
rect 26238 23042 26290 23054
rect 26238 22978 26290 22990
rect 27694 23042 27746 23054
rect 38558 23042 38610 23054
rect 28690 22990 28702 23042
rect 28754 22990 28766 23042
rect 31154 22990 31166 23042
rect 31218 22990 31230 23042
rect 27694 22978 27746 22990
rect 38558 22978 38610 22990
rect 16270 22930 16322 22942
rect 16270 22866 16322 22878
rect 21646 22930 21698 22942
rect 21646 22866 21698 22878
rect 25902 22930 25954 22942
rect 25902 22866 25954 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 9998 22594 10050 22606
rect 9998 22530 10050 22542
rect 28590 22594 28642 22606
rect 28590 22530 28642 22542
rect 29486 22594 29538 22606
rect 29486 22530 29538 22542
rect 29710 22594 29762 22606
rect 29710 22530 29762 22542
rect 29934 22594 29986 22606
rect 29934 22530 29986 22542
rect 34414 22594 34466 22606
rect 34414 22530 34466 22542
rect 4846 22482 4898 22494
rect 4846 22418 4898 22430
rect 5742 22482 5794 22494
rect 5742 22418 5794 22430
rect 6750 22482 6802 22494
rect 7534 22482 7586 22494
rect 8654 22482 8706 22494
rect 7186 22430 7198 22482
rect 7250 22430 7262 22482
rect 7970 22430 7982 22482
rect 8034 22430 8046 22482
rect 6750 22418 6802 22430
rect 7534 22418 7586 22430
rect 8654 22418 8706 22430
rect 11454 22482 11506 22494
rect 21646 22482 21698 22494
rect 25678 22482 25730 22494
rect 16146 22430 16158 22482
rect 16210 22430 16222 22482
rect 17378 22430 17390 22482
rect 17442 22430 17454 22482
rect 22194 22430 22206 22482
rect 22258 22430 22270 22482
rect 23090 22430 23102 22482
rect 23154 22430 23166 22482
rect 11454 22418 11506 22430
rect 21646 22418 21698 22430
rect 25678 22418 25730 22430
rect 27134 22482 27186 22494
rect 27134 22418 27186 22430
rect 27918 22482 27970 22494
rect 27918 22418 27970 22430
rect 30158 22482 30210 22494
rect 30158 22418 30210 22430
rect 30606 22482 30658 22494
rect 30606 22418 30658 22430
rect 31614 22482 31666 22494
rect 31614 22418 31666 22430
rect 35870 22482 35922 22494
rect 40002 22430 40014 22482
rect 40066 22430 40078 22482
rect 35870 22418 35922 22430
rect 3838 22370 3890 22382
rect 2818 22318 2830 22370
rect 2882 22318 2894 22370
rect 3838 22306 3890 22318
rect 8318 22370 8370 22382
rect 8318 22306 8370 22318
rect 9214 22370 9266 22382
rect 9214 22306 9266 22318
rect 11230 22370 11282 22382
rect 17054 22370 17106 22382
rect 18062 22370 18114 22382
rect 25790 22370 25842 22382
rect 29038 22370 29090 22382
rect 12002 22318 12014 22370
rect 12066 22318 12078 22370
rect 12674 22318 12686 22370
rect 12738 22318 12750 22370
rect 15922 22318 15934 22370
rect 15986 22318 15998 22370
rect 17602 22318 17614 22370
rect 17666 22318 17678 22370
rect 23314 22318 23326 22370
rect 23378 22318 23390 22370
rect 26226 22318 26238 22370
rect 26290 22318 26302 22370
rect 11230 22306 11282 22318
rect 17054 22306 17106 22318
rect 18062 22306 18114 22318
rect 25790 22306 25842 22318
rect 29038 22306 29090 22318
rect 32958 22370 33010 22382
rect 32958 22306 33010 22318
rect 33182 22370 33234 22382
rect 33182 22306 33234 22318
rect 34974 22370 35026 22382
rect 39106 22318 39118 22370
rect 39170 22318 39182 22370
rect 34974 22306 35026 22318
rect 1934 22258 1986 22270
rect 1934 22194 1986 22206
rect 3278 22258 3330 22270
rect 3278 22194 3330 22206
rect 6190 22258 6242 22270
rect 6190 22194 6242 22206
rect 8094 22258 8146 22270
rect 8094 22194 8146 22206
rect 9550 22258 9602 22270
rect 9550 22194 9602 22206
rect 9886 22258 9938 22270
rect 16606 22258 16658 22270
rect 12898 22206 12910 22258
rect 12962 22206 12974 22258
rect 9886 22194 9938 22206
rect 16606 22194 16658 22206
rect 17166 22258 17218 22270
rect 17166 22194 17218 22206
rect 18622 22258 18674 22270
rect 18622 22194 18674 22206
rect 21758 22258 21810 22270
rect 21758 22194 21810 22206
rect 22430 22258 22482 22270
rect 22430 22194 22482 22206
rect 28478 22258 28530 22270
rect 28478 22194 28530 22206
rect 32286 22258 32338 22270
rect 32286 22194 32338 22206
rect 33406 22258 33458 22270
rect 33406 22194 33458 22206
rect 33854 22258 33906 22270
rect 33854 22194 33906 22206
rect 33966 22258 34018 22270
rect 33966 22194 34018 22206
rect 34526 22258 34578 22270
rect 34526 22194 34578 22206
rect 35422 22258 35474 22270
rect 35422 22194 35474 22206
rect 2158 22146 2210 22158
rect 2158 22082 2210 22094
rect 4734 22146 4786 22158
rect 4734 22082 4786 22094
rect 6302 22146 6354 22158
rect 6302 22082 6354 22094
rect 7310 22146 7362 22158
rect 7310 22082 7362 22094
rect 8766 22146 8818 22158
rect 8766 22082 8818 22094
rect 8878 22146 8930 22158
rect 8878 22082 8930 22094
rect 9438 22146 9490 22158
rect 9438 22082 9490 22094
rect 10446 22146 10498 22158
rect 14142 22146 14194 22158
rect 10882 22094 10894 22146
rect 10946 22094 10958 22146
rect 11890 22094 11902 22146
rect 11954 22094 11966 22146
rect 10446 22082 10498 22094
rect 14142 22082 14194 22094
rect 14590 22146 14642 22158
rect 14590 22082 14642 22094
rect 17390 22146 17442 22158
rect 17390 22082 17442 22094
rect 18174 22146 18226 22158
rect 18174 22082 18226 22094
rect 18398 22146 18450 22158
rect 18398 22082 18450 22094
rect 18734 22146 18786 22158
rect 18734 22082 18786 22094
rect 18958 22146 19010 22158
rect 18958 22082 19010 22094
rect 19294 22146 19346 22158
rect 19294 22082 19346 22094
rect 19742 22146 19794 22158
rect 19742 22082 19794 22094
rect 20302 22146 20354 22158
rect 20302 22082 20354 22094
rect 20750 22146 20802 22158
rect 20750 22082 20802 22094
rect 21534 22146 21586 22158
rect 21534 22082 21586 22094
rect 22206 22146 22258 22158
rect 22206 22082 22258 22094
rect 27470 22146 27522 22158
rect 27470 22082 27522 22094
rect 31054 22146 31106 22158
rect 31054 22082 31106 22094
rect 33294 22146 33346 22158
rect 33294 22082 33346 22094
rect 33630 22146 33682 22158
rect 33630 22082 33682 22094
rect 34414 22146 34466 22158
rect 34414 22082 34466 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 1598 21810 1650 21822
rect 5630 21810 5682 21822
rect 2370 21758 2382 21810
rect 2434 21758 2446 21810
rect 1598 21746 1650 21758
rect 5630 21746 5682 21758
rect 8542 21810 8594 21822
rect 8542 21746 8594 21758
rect 9550 21810 9602 21822
rect 14702 21810 14754 21822
rect 12898 21758 12910 21810
rect 12962 21758 12974 21810
rect 13682 21758 13694 21810
rect 13746 21758 13758 21810
rect 9550 21746 9602 21758
rect 14702 21746 14754 21758
rect 17502 21810 17554 21822
rect 17502 21746 17554 21758
rect 17614 21810 17666 21822
rect 17614 21746 17666 21758
rect 25342 21810 25394 21822
rect 25342 21746 25394 21758
rect 30942 21810 30994 21822
rect 30942 21746 30994 21758
rect 33742 21810 33794 21822
rect 38222 21810 38274 21822
rect 37426 21758 37438 21810
rect 37490 21758 37502 21810
rect 33742 21746 33794 21758
rect 38222 21746 38274 21758
rect 5742 21698 5794 21710
rect 8766 21698 8818 21710
rect 14478 21698 14530 21710
rect 7746 21646 7758 21698
rect 7810 21646 7822 21698
rect 10098 21646 10110 21698
rect 10162 21646 10174 21698
rect 10434 21646 10446 21698
rect 10498 21646 10510 21698
rect 12562 21646 12574 21698
rect 12626 21646 12638 21698
rect 5742 21634 5794 21646
rect 8766 21634 8818 21646
rect 14478 21634 14530 21646
rect 15822 21698 15874 21710
rect 15822 21634 15874 21646
rect 24222 21698 24274 21710
rect 27918 21698 27970 21710
rect 27570 21646 27582 21698
rect 27634 21646 27646 21698
rect 24222 21634 24274 21646
rect 27918 21634 27970 21646
rect 29262 21698 29314 21710
rect 29262 21634 29314 21646
rect 32174 21698 32226 21710
rect 32174 21634 32226 21646
rect 33854 21698 33906 21710
rect 33854 21634 33906 21646
rect 38334 21698 38386 21710
rect 38334 21634 38386 21646
rect 5294 21586 5346 21598
rect 4722 21534 4734 21586
rect 4786 21534 4798 21586
rect 5294 21522 5346 21534
rect 5406 21586 5458 21598
rect 8318 21586 8370 21598
rect 6178 21534 6190 21586
rect 6242 21534 6254 21586
rect 6514 21534 6526 21586
rect 6578 21534 6590 21586
rect 8082 21534 8094 21586
rect 8146 21534 8158 21586
rect 5406 21522 5458 21534
rect 8318 21522 8370 21534
rect 9774 21586 9826 21598
rect 14366 21586 14418 21598
rect 12338 21534 12350 21586
rect 12402 21534 12414 21586
rect 13458 21534 13470 21586
rect 13522 21534 13534 21586
rect 9774 21522 9826 21534
rect 14366 21522 14418 21534
rect 15262 21586 15314 21598
rect 15262 21522 15314 21534
rect 15934 21586 15986 21598
rect 24334 21586 24386 21598
rect 30158 21586 30210 21598
rect 16482 21534 16494 21586
rect 16546 21534 16558 21586
rect 18498 21534 18510 21586
rect 18562 21534 18574 21586
rect 25666 21534 25678 21586
rect 25730 21534 25742 21586
rect 26898 21534 26910 21586
rect 26962 21534 26974 21586
rect 28354 21534 28366 21586
rect 28418 21534 28430 21586
rect 29698 21534 29710 21586
rect 29762 21534 29774 21586
rect 15934 21522 15986 21534
rect 24334 21522 24386 21534
rect 30158 21522 30210 21534
rect 30606 21586 30658 21598
rect 30606 21522 30658 21534
rect 30830 21586 30882 21598
rect 30830 21522 30882 21534
rect 31166 21586 31218 21598
rect 33966 21586 34018 21598
rect 32498 21534 32510 21586
rect 32562 21534 32574 21586
rect 33618 21534 33630 21586
rect 33682 21534 33694 21586
rect 31166 21522 31218 21534
rect 33966 21522 34018 21534
rect 34526 21586 34578 21598
rect 34850 21534 34862 21586
rect 34914 21534 34926 21586
rect 38994 21534 39006 21586
rect 39058 21534 39070 21586
rect 34526 21522 34578 21534
rect 10558 21474 10610 21486
rect 8194 21422 8206 21474
rect 8258 21422 8270 21474
rect 10558 21410 10610 21422
rect 11006 21474 11058 21486
rect 11006 21410 11058 21422
rect 15486 21474 15538 21486
rect 15486 21410 15538 21422
rect 18286 21474 18338 21486
rect 31726 21474 31778 21486
rect 22306 21422 22318 21474
rect 22370 21422 22382 21474
rect 28802 21422 28814 21474
rect 28866 21422 28878 21474
rect 40114 21422 40126 21474
rect 40178 21422 40190 21474
rect 18286 21410 18338 21422
rect 31726 21410 31778 21422
rect 17726 21362 17778 21374
rect 14914 21310 14926 21362
rect 14978 21310 14990 21362
rect 17726 21298 17778 21310
rect 24222 21362 24274 21374
rect 24222 21298 24274 21310
rect 31838 21362 31890 21374
rect 31838 21298 31890 21310
rect 32510 21362 32562 21374
rect 32510 21298 32562 21310
rect 33070 21362 33122 21374
rect 33070 21298 33122 21310
rect 33294 21362 33346 21374
rect 33294 21298 33346 21310
rect 37998 21362 38050 21374
rect 37998 21298 38050 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 11790 21026 11842 21038
rect 14478 21026 14530 21038
rect 20638 21026 20690 21038
rect 12674 20974 12686 21026
rect 12738 20974 12750 21026
rect 19058 20974 19070 21026
rect 19122 21023 19134 21026
rect 19618 21023 19630 21026
rect 19122 20977 19630 21023
rect 19122 20974 19134 20977
rect 19618 20974 19630 20977
rect 19682 20974 19694 21026
rect 11790 20962 11842 20974
rect 14478 20962 14530 20974
rect 20638 20962 20690 20974
rect 27582 21026 27634 21038
rect 27582 20962 27634 20974
rect 29262 21026 29314 21038
rect 33070 21026 33122 21038
rect 35422 21026 35474 21038
rect 31490 20974 31502 21026
rect 31554 20974 31566 21026
rect 33954 20974 33966 21026
rect 34018 20974 34030 21026
rect 29262 20962 29314 20974
rect 33070 20962 33122 20974
rect 35422 20962 35474 20974
rect 3726 20914 3778 20926
rect 3726 20850 3778 20862
rect 4622 20914 4674 20926
rect 4622 20850 4674 20862
rect 6302 20914 6354 20926
rect 6302 20850 6354 20862
rect 7982 20914 8034 20926
rect 19294 20914 19346 20926
rect 18610 20862 18622 20914
rect 18674 20862 18686 20914
rect 7982 20850 8034 20862
rect 19294 20850 19346 20862
rect 20190 20914 20242 20926
rect 20190 20850 20242 20862
rect 22878 20914 22930 20926
rect 22878 20850 22930 20862
rect 24222 20914 24274 20926
rect 26686 20914 26738 20926
rect 24658 20862 24670 20914
rect 24722 20862 24734 20914
rect 25442 20862 25454 20914
rect 25506 20862 25518 20914
rect 24222 20850 24274 20862
rect 26686 20850 26738 20862
rect 29822 20914 29874 20926
rect 29822 20850 29874 20862
rect 30942 20914 30994 20926
rect 30942 20850 30994 20862
rect 31950 20914 32002 20926
rect 31950 20850 32002 20862
rect 33630 20914 33682 20926
rect 33630 20850 33682 20862
rect 35534 20914 35586 20926
rect 35534 20850 35586 20862
rect 1710 20802 1762 20814
rect 1710 20738 1762 20750
rect 4286 20802 4338 20814
rect 4286 20738 4338 20750
rect 4510 20802 4562 20814
rect 4510 20738 4562 20750
rect 5182 20802 5234 20814
rect 5182 20738 5234 20750
rect 6190 20802 6242 20814
rect 6974 20802 7026 20814
rect 8878 20802 8930 20814
rect 6738 20750 6750 20802
rect 6802 20750 6814 20802
rect 8418 20750 8430 20802
rect 8482 20750 8494 20802
rect 6190 20738 6242 20750
rect 6974 20738 7026 20750
rect 8878 20738 8930 20750
rect 9662 20802 9714 20814
rect 9662 20738 9714 20750
rect 12126 20802 12178 20814
rect 12126 20738 12178 20750
rect 12350 20802 12402 20814
rect 12350 20738 12402 20750
rect 13470 20802 13522 20814
rect 13470 20738 13522 20750
rect 13694 20802 13746 20814
rect 13694 20738 13746 20750
rect 13918 20802 13970 20814
rect 15710 20802 15762 20814
rect 17054 20802 17106 20814
rect 15362 20750 15374 20802
rect 15426 20750 15438 20802
rect 16482 20750 16494 20802
rect 16546 20750 16558 20802
rect 13918 20738 13970 20750
rect 15710 20738 15762 20750
rect 17054 20738 17106 20750
rect 17614 20802 17666 20814
rect 17614 20738 17666 20750
rect 18062 20802 18114 20814
rect 18062 20738 18114 20750
rect 20750 20802 20802 20814
rect 20750 20738 20802 20750
rect 22654 20802 22706 20814
rect 22654 20738 22706 20750
rect 23102 20802 23154 20814
rect 23102 20738 23154 20750
rect 23326 20802 23378 20814
rect 23326 20738 23378 20750
rect 23998 20802 24050 20814
rect 31166 20802 31218 20814
rect 25778 20750 25790 20802
rect 25842 20750 25854 20802
rect 27682 20750 27694 20802
rect 27746 20750 27758 20802
rect 23998 20738 24050 20750
rect 31166 20738 31218 20750
rect 32846 20802 32898 20814
rect 35086 20802 35138 20814
rect 33730 20750 33742 20802
rect 33794 20750 33806 20802
rect 34402 20750 34414 20802
rect 34466 20750 34478 20802
rect 32846 20738 32898 20750
rect 35086 20738 35138 20750
rect 35198 20802 35250 20814
rect 35198 20738 35250 20750
rect 37886 20802 37938 20814
rect 37886 20738 37938 20750
rect 2270 20690 2322 20702
rect 2270 20626 2322 20638
rect 3166 20690 3218 20702
rect 3166 20626 3218 20638
rect 4734 20690 4786 20702
rect 4734 20626 4786 20638
rect 7422 20690 7474 20702
rect 7422 20626 7474 20638
rect 9550 20690 9602 20702
rect 11678 20690 11730 20702
rect 10210 20638 10222 20690
rect 10274 20638 10286 20690
rect 10434 20638 10446 20690
rect 10498 20638 10510 20690
rect 9550 20626 9602 20638
rect 11678 20626 11730 20638
rect 14366 20690 14418 20702
rect 14366 20626 14418 20638
rect 15822 20690 15874 20702
rect 15822 20626 15874 20638
rect 17166 20690 17218 20702
rect 17166 20626 17218 20638
rect 18846 20690 18898 20702
rect 18846 20626 18898 20638
rect 19854 20690 19906 20702
rect 19854 20626 19906 20638
rect 20638 20690 20690 20702
rect 20638 20626 20690 20638
rect 21758 20690 21810 20702
rect 29150 20690 29202 20702
rect 22082 20638 22094 20690
rect 22146 20638 22158 20690
rect 27346 20638 27358 20690
rect 27410 20638 27422 20690
rect 21758 20626 21810 20638
rect 29150 20626 29202 20638
rect 40238 20690 40290 20702
rect 40238 20626 40290 20638
rect 2606 20578 2658 20590
rect 2606 20514 2658 20526
rect 5966 20578 6018 20590
rect 5966 20514 6018 20526
rect 6414 20578 6466 20590
rect 6414 20514 6466 20526
rect 7534 20578 7586 20590
rect 7534 20514 7586 20526
rect 7646 20578 7698 20590
rect 7646 20514 7698 20526
rect 13582 20578 13634 20590
rect 13582 20514 13634 20526
rect 17726 20578 17778 20590
rect 17726 20514 17778 20526
rect 17838 20578 17890 20590
rect 17838 20514 17890 20526
rect 17950 20578 18002 20590
rect 17950 20514 18002 20526
rect 18622 20578 18674 20590
rect 18622 20514 18674 20526
rect 21422 20578 21474 20590
rect 28142 20578 28194 20590
rect 23650 20526 23662 20578
rect 23714 20526 23726 20578
rect 21422 20514 21474 20526
rect 28142 20514 28194 20526
rect 28590 20578 28642 20590
rect 28590 20514 28642 20526
rect 29262 20578 29314 20590
rect 29262 20514 29314 20526
rect 30270 20578 30322 20590
rect 30270 20514 30322 20526
rect 32398 20578 32450 20590
rect 32398 20514 32450 20526
rect 32510 20578 32562 20590
rect 32510 20514 32562 20526
rect 32622 20578 32674 20590
rect 32622 20514 32674 20526
rect 36094 20578 36146 20590
rect 36094 20514 36146 20526
rect 39678 20578 39730 20590
rect 39678 20514 39730 20526
rect 39902 20578 39954 20590
rect 39902 20514 39954 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 4734 20242 4786 20254
rect 4734 20178 4786 20190
rect 5742 20242 5794 20254
rect 5742 20178 5794 20190
rect 9662 20242 9714 20254
rect 9662 20178 9714 20190
rect 10334 20242 10386 20254
rect 17726 20242 17778 20254
rect 14018 20190 14030 20242
rect 14082 20190 14094 20242
rect 10334 20178 10386 20190
rect 17726 20178 17778 20190
rect 17838 20242 17890 20254
rect 17838 20178 17890 20190
rect 18622 20242 18674 20254
rect 24446 20242 24498 20254
rect 30606 20242 30658 20254
rect 23426 20190 23438 20242
rect 23490 20190 23502 20242
rect 25218 20190 25230 20242
rect 25282 20190 25294 20242
rect 18622 20178 18674 20190
rect 24446 20178 24498 20190
rect 30606 20178 30658 20190
rect 3614 20130 3666 20142
rect 3614 20066 3666 20078
rect 5182 20130 5234 20142
rect 5182 20066 5234 20078
rect 5630 20130 5682 20142
rect 5630 20066 5682 20078
rect 6414 20130 6466 20142
rect 6414 20066 6466 20078
rect 8206 20130 8258 20142
rect 8206 20066 8258 20078
rect 9774 20130 9826 20142
rect 9774 20066 9826 20078
rect 14142 20130 14194 20142
rect 18062 20130 18114 20142
rect 16706 20078 16718 20130
rect 16770 20078 16782 20130
rect 14142 20066 14194 20078
rect 18062 20066 18114 20078
rect 24222 20130 24274 20142
rect 24222 20066 24274 20078
rect 26238 20130 26290 20142
rect 37662 20130 37714 20142
rect 29138 20078 29150 20130
rect 29202 20078 29214 20130
rect 33394 20078 33406 20130
rect 33458 20078 33470 20130
rect 26238 20066 26290 20078
rect 37662 20066 37714 20078
rect 38446 20130 38498 20142
rect 38446 20066 38498 20078
rect 7870 20018 7922 20030
rect 2706 19966 2718 20018
rect 2770 19966 2782 20018
rect 6178 19966 6190 20018
rect 6242 19966 6254 20018
rect 7298 19966 7310 20018
rect 7362 19966 7374 20018
rect 7870 19954 7922 19966
rect 8430 20018 8482 20030
rect 8430 19954 8482 19966
rect 8654 20018 8706 20030
rect 10446 20018 10498 20030
rect 8866 19966 8878 20018
rect 8930 19966 8942 20018
rect 8654 19954 8706 19966
rect 10446 19954 10498 19966
rect 14702 20018 14754 20030
rect 17614 20018 17666 20030
rect 20526 20018 20578 20030
rect 24782 20018 24834 20030
rect 15026 19966 15038 20018
rect 15090 19966 15102 20018
rect 17378 19966 17390 20018
rect 17442 19966 17454 20018
rect 19842 19966 19854 20018
rect 19906 19966 19918 20018
rect 20962 19966 20974 20018
rect 21026 19966 21038 20018
rect 14702 19954 14754 19966
rect 17614 19954 17666 19966
rect 20526 19954 20578 19966
rect 24782 19954 24834 19966
rect 25566 20018 25618 20030
rect 25566 19954 25618 19966
rect 26574 20018 26626 20030
rect 26574 19954 26626 19966
rect 26686 20018 26738 20030
rect 26686 19954 26738 19966
rect 26798 20018 26850 20030
rect 26798 19954 26850 19966
rect 27246 20018 27298 20030
rect 27246 19954 27298 19966
rect 30382 20018 30434 20030
rect 30382 19954 30434 19966
rect 31950 20018 32002 20030
rect 34078 20018 34130 20030
rect 33618 19966 33630 20018
rect 33682 19966 33694 20018
rect 31950 19954 32002 19966
rect 34078 19954 34130 19966
rect 34974 20018 35026 20030
rect 35298 19966 35310 20018
rect 35362 19966 35374 20018
rect 38994 19966 39006 20018
rect 39058 19966 39070 20018
rect 34974 19954 35026 19966
rect 4062 19906 4114 19918
rect 1922 19854 1934 19906
rect 1986 19854 1998 19906
rect 4062 19842 4114 19854
rect 6526 19906 6578 19918
rect 9550 19906 9602 19918
rect 7074 19854 7086 19906
rect 7138 19854 7150 19906
rect 8754 19854 8766 19906
rect 8818 19854 8830 19906
rect 6526 19842 6578 19854
rect 9550 19842 9602 19854
rect 10894 19906 10946 19918
rect 10894 19842 10946 19854
rect 12238 19906 12290 19918
rect 12238 19842 12290 19854
rect 12686 19906 12738 19918
rect 25790 19906 25842 19918
rect 19170 19854 19182 19906
rect 19234 19854 19246 19906
rect 12686 19842 12738 19854
rect 25790 19842 25842 19854
rect 27582 19906 27634 19918
rect 27582 19842 27634 19854
rect 28030 19906 28082 19918
rect 28030 19842 28082 19854
rect 28478 19906 28530 19918
rect 28478 19842 28530 19854
rect 31502 19906 31554 19918
rect 31502 19842 31554 19854
rect 32510 19906 32562 19918
rect 40002 19854 40014 19906
rect 40066 19854 40078 19906
rect 32510 19842 32562 19854
rect 5854 19794 5906 19806
rect 5854 19730 5906 19742
rect 10334 19794 10386 19806
rect 10334 19730 10386 19742
rect 23998 19794 24050 19806
rect 23998 19730 24050 19742
rect 24558 19794 24610 19806
rect 24558 19730 24610 19742
rect 26126 19794 26178 19806
rect 26126 19730 26178 19742
rect 29710 19794 29762 19806
rect 29710 19730 29762 19742
rect 29934 19794 29986 19806
rect 29934 19730 29986 19742
rect 30158 19794 30210 19806
rect 30158 19730 30210 19742
rect 31054 19794 31106 19806
rect 31054 19730 31106 19742
rect 31278 19794 31330 19806
rect 31278 19730 31330 19742
rect 34414 19794 34466 19806
rect 34414 19730 34466 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 8542 19458 8594 19470
rect 12798 19458 12850 19470
rect 8866 19406 8878 19458
rect 8930 19406 8942 19458
rect 8542 19394 8594 19406
rect 12798 19394 12850 19406
rect 14254 19458 14306 19470
rect 14254 19394 14306 19406
rect 14478 19458 14530 19470
rect 14478 19394 14530 19406
rect 20862 19458 20914 19470
rect 20862 19394 20914 19406
rect 23774 19458 23826 19470
rect 23774 19394 23826 19406
rect 25342 19458 25394 19470
rect 25342 19394 25394 19406
rect 25678 19458 25730 19470
rect 37662 19458 37714 19470
rect 34290 19406 34302 19458
rect 34354 19406 34366 19458
rect 25678 19394 25730 19406
rect 37662 19394 37714 19406
rect 4174 19346 4226 19358
rect 8318 19346 8370 19358
rect 7746 19294 7758 19346
rect 7810 19294 7822 19346
rect 4174 19282 4226 19294
rect 8318 19282 8370 19294
rect 11566 19346 11618 19358
rect 15934 19346 15986 19358
rect 31166 19346 31218 19358
rect 35534 19346 35586 19358
rect 15138 19294 15150 19346
rect 15202 19294 15214 19346
rect 22194 19294 22206 19346
rect 22258 19294 22270 19346
rect 30258 19294 30270 19346
rect 30322 19294 30334 19346
rect 34178 19294 34190 19346
rect 34242 19294 34254 19346
rect 11566 19282 11618 19294
rect 15934 19282 15986 19294
rect 31166 19282 31218 19294
rect 35534 19282 35586 19294
rect 37214 19346 37266 19358
rect 37214 19282 37266 19294
rect 37550 19346 37602 19358
rect 37550 19282 37602 19294
rect 4510 19234 4562 19246
rect 2930 19182 2942 19234
rect 2994 19182 3006 19234
rect 3378 19182 3390 19234
rect 3442 19182 3454 19234
rect 4510 19170 4562 19182
rect 4734 19234 4786 19246
rect 4734 19170 4786 19182
rect 5182 19234 5234 19246
rect 5182 19170 5234 19182
rect 5518 19234 5570 19246
rect 5518 19170 5570 19182
rect 5854 19234 5906 19246
rect 11678 19234 11730 19246
rect 6290 19182 6302 19234
rect 6354 19182 6366 19234
rect 6850 19182 6862 19234
rect 6914 19182 6926 19234
rect 10994 19182 11006 19234
rect 11058 19182 11070 19234
rect 5854 19170 5906 19182
rect 11678 19170 11730 19182
rect 11902 19234 11954 19246
rect 12462 19234 12514 19246
rect 12114 19182 12126 19234
rect 12178 19182 12190 19234
rect 11902 19170 11954 19182
rect 12462 19170 12514 19182
rect 12910 19234 12962 19246
rect 16718 19234 16770 19246
rect 15250 19182 15262 19234
rect 15314 19182 15326 19234
rect 12910 19170 12962 19182
rect 16718 19170 16770 19182
rect 16830 19234 16882 19246
rect 16830 19170 16882 19182
rect 16942 19234 16994 19246
rect 16942 19170 16994 19182
rect 17166 19234 17218 19246
rect 24110 19234 24162 19246
rect 26126 19234 26178 19246
rect 17714 19182 17726 19234
rect 17778 19182 17790 19234
rect 23090 19182 23102 19234
rect 23154 19182 23166 19234
rect 24658 19182 24670 19234
rect 24722 19182 24734 19234
rect 25666 19182 25678 19234
rect 25730 19182 25742 19234
rect 17166 19170 17218 19182
rect 24110 19170 24162 19182
rect 26126 19170 26178 19182
rect 26350 19234 26402 19246
rect 30718 19234 30770 19246
rect 34750 19234 34802 19246
rect 28466 19182 28478 19234
rect 28530 19182 28542 19234
rect 33730 19182 33742 19234
rect 33794 19182 33806 19234
rect 26350 19170 26402 19182
rect 30718 19170 30770 19182
rect 34750 19170 34802 19182
rect 5742 19122 5794 19134
rect 11454 19122 11506 19134
rect 2034 19070 2046 19122
rect 2098 19070 2110 19122
rect 3602 19070 3614 19122
rect 3666 19070 3678 19122
rect 10770 19070 10782 19122
rect 10834 19070 10846 19122
rect 5742 19058 5794 19070
rect 11454 19058 11506 19070
rect 13694 19122 13746 19134
rect 13694 19058 13746 19070
rect 13918 19122 13970 19134
rect 13918 19058 13970 19070
rect 14030 19122 14082 19134
rect 14030 19058 14082 19070
rect 21422 19122 21474 19134
rect 26238 19122 26290 19134
rect 24882 19070 24894 19122
rect 24946 19070 24958 19122
rect 21422 19058 21474 19070
rect 26238 19058 26290 19070
rect 26574 19122 26626 19134
rect 26574 19058 26626 19070
rect 31054 19122 31106 19134
rect 31054 19058 31106 19070
rect 32622 19122 32674 19134
rect 32622 19058 32674 19070
rect 35086 19122 35138 19134
rect 35086 19058 35138 19070
rect 40238 19122 40290 19134
rect 40238 19058 40290 19070
rect 4622 19010 4674 19022
rect 4622 18946 4674 18958
rect 9326 19010 9378 19022
rect 9326 18946 9378 18958
rect 9774 19010 9826 19022
rect 9774 18946 9826 18958
rect 10222 19010 10274 19022
rect 10222 18946 10274 18958
rect 12798 19010 12850 19022
rect 12798 18946 12850 18958
rect 16494 19010 16546 19022
rect 21310 19010 21362 19022
rect 20290 18958 20302 19010
rect 20354 18958 20366 19010
rect 16494 18946 16546 18958
rect 21310 18946 21362 18958
rect 28030 19010 28082 19022
rect 28030 18946 28082 18958
rect 29262 19010 29314 19022
rect 29262 18946 29314 18958
rect 31278 19010 31330 19022
rect 31278 18946 31330 18958
rect 31502 19010 31554 19022
rect 31502 18946 31554 18958
rect 32062 19010 32114 19022
rect 32062 18946 32114 18958
rect 32734 19010 32786 19022
rect 32734 18946 32786 18958
rect 35982 19010 36034 19022
rect 35982 18946 36034 18958
rect 39678 19010 39730 19022
rect 39678 18946 39730 18958
rect 39902 19010 39954 19022
rect 39902 18946 39954 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 5630 18674 5682 18686
rect 4946 18622 4958 18674
rect 5010 18622 5022 18674
rect 5630 18610 5682 18622
rect 6190 18674 6242 18686
rect 6190 18610 6242 18622
rect 7982 18674 8034 18686
rect 7982 18610 8034 18622
rect 8766 18674 8818 18686
rect 8766 18610 8818 18622
rect 13134 18674 13186 18686
rect 13134 18610 13186 18622
rect 13358 18674 13410 18686
rect 13358 18610 13410 18622
rect 15038 18674 15090 18686
rect 15038 18610 15090 18622
rect 15934 18674 15986 18686
rect 15934 18610 15986 18622
rect 17726 18674 17778 18686
rect 17726 18610 17778 18622
rect 18062 18674 18114 18686
rect 18062 18610 18114 18622
rect 18734 18674 18786 18686
rect 18734 18610 18786 18622
rect 24222 18674 24274 18686
rect 24222 18610 24274 18622
rect 24558 18674 24610 18686
rect 24558 18610 24610 18622
rect 6302 18562 6354 18574
rect 6302 18498 6354 18510
rect 6862 18562 6914 18574
rect 6862 18498 6914 18510
rect 6974 18562 7026 18574
rect 6974 18498 7026 18510
rect 7534 18562 7586 18574
rect 7534 18498 7586 18510
rect 8318 18562 8370 18574
rect 8318 18498 8370 18510
rect 12014 18562 12066 18574
rect 12014 18498 12066 18510
rect 14030 18562 14082 18574
rect 14030 18498 14082 18510
rect 14254 18562 14306 18574
rect 14254 18498 14306 18510
rect 14926 18562 14978 18574
rect 14926 18498 14978 18510
rect 15822 18562 15874 18574
rect 22866 18510 22878 18562
rect 22930 18510 22942 18562
rect 15822 18498 15874 18510
rect 2158 18450 2210 18462
rect 8542 18450 8594 18462
rect 9550 18450 9602 18462
rect 10446 18450 10498 18462
rect 13022 18450 13074 18462
rect 15262 18450 15314 18462
rect 2594 18398 2606 18450
rect 2658 18398 2670 18450
rect 8978 18398 8990 18450
rect 9042 18398 9054 18450
rect 10210 18398 10222 18450
rect 10274 18398 10286 18450
rect 11106 18398 11118 18450
rect 11170 18398 11182 18450
rect 13570 18398 13582 18450
rect 13634 18398 13646 18450
rect 2158 18386 2210 18398
rect 8542 18386 8594 18398
rect 9550 18386 9602 18398
rect 10446 18386 10498 18398
rect 13022 18386 13074 18398
rect 15262 18386 15314 18398
rect 15374 18450 15426 18462
rect 15374 18386 15426 18398
rect 16270 18450 16322 18462
rect 16270 18386 16322 18398
rect 17838 18450 17890 18462
rect 17838 18386 17890 18398
rect 18174 18450 18226 18462
rect 18174 18386 18226 18398
rect 19182 18450 19234 18462
rect 23214 18450 23266 18462
rect 19730 18398 19742 18450
rect 19794 18398 19806 18450
rect 21634 18398 21646 18450
rect 21698 18398 21710 18450
rect 19182 18386 19234 18398
rect 23214 18386 23266 18398
rect 23550 18450 23602 18462
rect 26910 18450 26962 18462
rect 25442 18398 25454 18450
rect 25506 18398 25518 18450
rect 23550 18386 23602 18398
rect 26910 18386 26962 18398
rect 33182 18450 33234 18462
rect 33842 18398 33854 18450
rect 33906 18398 33918 18450
rect 33182 18386 33234 18398
rect 12574 18338 12626 18350
rect 8866 18286 8878 18338
rect 8930 18286 8942 18338
rect 12114 18286 12126 18338
rect 12178 18286 12190 18338
rect 12574 18274 12626 18286
rect 13246 18338 13298 18350
rect 16382 18338 16434 18350
rect 13906 18286 13918 18338
rect 13970 18286 13982 18338
rect 13246 18274 13298 18286
rect 16382 18274 16434 18286
rect 16830 18338 16882 18350
rect 21422 18338 21474 18350
rect 21982 18338 22034 18350
rect 20402 18286 20414 18338
rect 20466 18286 20478 18338
rect 21746 18286 21758 18338
rect 21810 18286 21822 18338
rect 16830 18274 16882 18286
rect 21422 18274 21474 18286
rect 21982 18274 22034 18286
rect 22430 18338 22482 18350
rect 22430 18274 22482 18286
rect 23662 18338 23714 18350
rect 26798 18338 26850 18350
rect 25890 18286 25902 18338
rect 25954 18286 25966 18338
rect 23662 18274 23714 18286
rect 26798 18274 26850 18286
rect 27358 18338 27410 18350
rect 27358 18274 27410 18286
rect 27806 18338 27858 18350
rect 27806 18274 27858 18286
rect 28254 18338 28306 18350
rect 28254 18274 28306 18286
rect 28702 18338 28754 18350
rect 28702 18274 28754 18286
rect 29150 18338 29202 18350
rect 29150 18274 29202 18286
rect 29710 18338 29762 18350
rect 29710 18274 29762 18286
rect 30046 18338 30098 18350
rect 30046 18274 30098 18286
rect 30718 18338 30770 18350
rect 30718 18274 30770 18286
rect 31166 18338 31218 18350
rect 31166 18274 31218 18286
rect 31726 18338 31778 18350
rect 31726 18274 31778 18286
rect 32174 18338 32226 18350
rect 34638 18338 34690 18350
rect 34066 18286 34078 18338
rect 34130 18286 34142 18338
rect 32174 18274 32226 18286
rect 34638 18274 34690 18286
rect 35086 18338 35138 18350
rect 35086 18274 35138 18286
rect 35534 18338 35586 18350
rect 35534 18274 35586 18286
rect 6974 18226 7026 18238
rect 6974 18162 7026 18174
rect 11118 18226 11170 18238
rect 11118 18162 11170 18174
rect 11454 18226 11506 18238
rect 11454 18162 11506 18174
rect 11790 18226 11842 18238
rect 11790 18162 11842 18174
rect 12462 18226 12514 18238
rect 34526 18226 34578 18238
rect 23874 18174 23886 18226
rect 23938 18223 23950 18226
rect 24658 18223 24670 18226
rect 23938 18177 24670 18223
rect 23938 18174 23950 18177
rect 24658 18174 24670 18177
rect 24722 18174 24734 18226
rect 28018 18174 28030 18226
rect 28082 18223 28094 18226
rect 28802 18223 28814 18226
rect 28082 18177 28814 18223
rect 28082 18174 28094 18177
rect 28802 18174 28814 18177
rect 28866 18174 28878 18226
rect 31266 18174 31278 18226
rect 31330 18223 31342 18226
rect 32610 18223 32622 18226
rect 31330 18177 32622 18223
rect 31330 18174 31342 18177
rect 32610 18174 32622 18177
rect 32674 18174 32686 18226
rect 12462 18162 12514 18174
rect 34526 18162 34578 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 4958 17890 5010 17902
rect 4958 17826 5010 17838
rect 13470 17890 13522 17902
rect 13470 17826 13522 17838
rect 13806 17890 13858 17902
rect 20414 17890 20466 17902
rect 17490 17838 17502 17890
rect 17554 17887 17566 17890
rect 18162 17887 18174 17890
rect 17554 17841 18174 17887
rect 17554 17838 17566 17841
rect 18162 17838 18174 17841
rect 18226 17838 18238 17890
rect 28018 17838 28030 17890
rect 28082 17887 28094 17890
rect 28242 17887 28254 17890
rect 28082 17841 28254 17887
rect 28082 17838 28094 17841
rect 28242 17838 28254 17841
rect 28306 17838 28318 17890
rect 13806 17826 13858 17838
rect 20414 17826 20466 17838
rect 2270 17778 2322 17790
rect 2270 17714 2322 17726
rect 3166 17778 3218 17790
rect 3166 17714 3218 17726
rect 5070 17778 5122 17790
rect 5070 17714 5122 17726
rect 6190 17778 6242 17790
rect 6190 17714 6242 17726
rect 6526 17778 6578 17790
rect 11454 17778 11506 17790
rect 10658 17726 10670 17778
rect 10722 17726 10734 17778
rect 6526 17714 6578 17726
rect 11454 17714 11506 17726
rect 11902 17778 11954 17790
rect 11902 17714 11954 17726
rect 14142 17778 14194 17790
rect 14142 17714 14194 17726
rect 14254 17778 14306 17790
rect 14254 17714 14306 17726
rect 16270 17778 16322 17790
rect 16270 17714 16322 17726
rect 16606 17778 16658 17790
rect 16606 17714 16658 17726
rect 17054 17778 17106 17790
rect 17054 17714 17106 17726
rect 18062 17778 18114 17790
rect 18062 17714 18114 17726
rect 18398 17778 18450 17790
rect 18398 17714 18450 17726
rect 18958 17778 19010 17790
rect 28030 17778 28082 17790
rect 19954 17726 19966 17778
rect 20018 17726 20030 17778
rect 21858 17726 21870 17778
rect 21922 17726 21934 17778
rect 23202 17726 23214 17778
rect 23266 17726 23278 17778
rect 18958 17714 19010 17726
rect 28030 17714 28082 17726
rect 29374 17778 29426 17790
rect 29374 17714 29426 17726
rect 34638 17778 34690 17790
rect 34638 17714 34690 17726
rect 35982 17778 36034 17790
rect 40002 17726 40014 17778
rect 40066 17726 40078 17778
rect 35982 17714 36034 17726
rect 4734 17666 4786 17678
rect 4734 17602 4786 17614
rect 8878 17666 8930 17678
rect 8878 17602 8930 17614
rect 9550 17666 9602 17678
rect 9550 17602 9602 17614
rect 9774 17666 9826 17678
rect 11790 17666 11842 17678
rect 10770 17614 10782 17666
rect 10834 17614 10846 17666
rect 9774 17602 9826 17614
rect 11790 17602 11842 17614
rect 12126 17666 12178 17678
rect 12126 17602 12178 17614
rect 12238 17666 12290 17678
rect 21310 17666 21362 17678
rect 23998 17666 24050 17678
rect 29710 17666 29762 17678
rect 33854 17666 33906 17678
rect 12562 17614 12574 17666
rect 12626 17614 12638 17666
rect 19842 17614 19854 17666
rect 19906 17614 19918 17666
rect 20290 17614 20302 17666
rect 20354 17614 20366 17666
rect 22754 17614 22766 17666
rect 22818 17614 22830 17666
rect 24658 17614 24670 17666
rect 24722 17614 24734 17666
rect 30370 17614 30382 17666
rect 30434 17614 30446 17666
rect 12238 17602 12290 17614
rect 21310 17602 21362 17614
rect 23998 17602 24050 17614
rect 29710 17602 29762 17614
rect 33854 17602 33906 17614
rect 34302 17666 34354 17678
rect 39106 17614 39118 17666
rect 39170 17614 39182 17666
rect 34302 17602 34354 17614
rect 1710 17554 1762 17566
rect 1710 17490 1762 17502
rect 3726 17554 3778 17566
rect 3726 17490 3778 17502
rect 10110 17554 10162 17566
rect 10110 17490 10162 17502
rect 14366 17554 14418 17566
rect 14366 17490 14418 17502
rect 14926 17554 14978 17566
rect 14926 17490 14978 17502
rect 35534 17554 35586 17566
rect 35534 17490 35586 17502
rect 2606 17442 2658 17454
rect 2606 17378 2658 17390
rect 4062 17442 4114 17454
rect 4062 17378 4114 17390
rect 8542 17442 8594 17454
rect 8542 17378 8594 17390
rect 8990 17442 9042 17454
rect 8990 17378 9042 17390
rect 9102 17442 9154 17454
rect 9102 17378 9154 17390
rect 9998 17442 10050 17454
rect 9998 17378 10050 17390
rect 13582 17442 13634 17454
rect 13582 17378 13634 17390
rect 15374 17442 15426 17454
rect 15374 17378 15426 17390
rect 17502 17442 17554 17454
rect 27694 17442 27746 17454
rect 26898 17390 26910 17442
rect 26962 17390 26974 17442
rect 17502 17378 17554 17390
rect 27694 17378 27746 17390
rect 28478 17442 28530 17454
rect 28478 17378 28530 17390
rect 29486 17442 29538 17454
rect 33406 17442 33458 17454
rect 32834 17390 32846 17442
rect 32898 17390 32910 17442
rect 29486 17378 29538 17390
rect 33406 17378 33458 17390
rect 33630 17442 33682 17454
rect 33630 17378 33682 17390
rect 33742 17442 33794 17454
rect 33742 17378 33794 17390
rect 34526 17442 34578 17454
rect 34526 17378 34578 17390
rect 35086 17442 35138 17454
rect 35086 17378 35138 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 1822 17106 1874 17118
rect 1822 17042 1874 17054
rect 2942 17106 2994 17118
rect 2942 17042 2994 17054
rect 10110 17106 10162 17118
rect 10110 17042 10162 17054
rect 12014 17106 12066 17118
rect 12014 17042 12066 17054
rect 14142 17106 14194 17118
rect 14142 17042 14194 17054
rect 15486 17106 15538 17118
rect 15486 17042 15538 17054
rect 19294 17106 19346 17118
rect 19294 17042 19346 17054
rect 23774 17106 23826 17118
rect 23774 17042 23826 17054
rect 24110 17106 24162 17118
rect 24110 17042 24162 17054
rect 26910 17106 26962 17118
rect 26910 17042 26962 17054
rect 33182 17106 33234 17118
rect 33182 17042 33234 17054
rect 10334 16994 10386 17006
rect 10334 16930 10386 16942
rect 11790 16994 11842 17006
rect 11790 16930 11842 16942
rect 12686 16994 12738 17006
rect 12686 16930 12738 16942
rect 14254 16994 14306 17006
rect 14254 16930 14306 16942
rect 14814 16994 14866 17006
rect 14814 16930 14866 16942
rect 17502 16994 17554 17006
rect 21086 16994 21138 17006
rect 24558 16994 24610 17006
rect 18386 16942 18398 16994
rect 18450 16942 18462 16994
rect 23090 16942 23102 16994
rect 23154 16942 23166 16994
rect 17502 16930 17554 16942
rect 21086 16930 21138 16942
rect 24558 16930 24610 16942
rect 33294 16994 33346 17006
rect 33294 16930 33346 16942
rect 36430 16994 36482 17006
rect 36430 16930 36482 16942
rect 37214 16994 37266 17006
rect 37214 16930 37266 16942
rect 12462 16882 12514 16894
rect 10994 16830 11006 16882
rect 11058 16830 11070 16882
rect 12462 16818 12514 16830
rect 12798 16882 12850 16894
rect 13918 16882 13970 16894
rect 13346 16830 13358 16882
rect 13410 16830 13422 16882
rect 12798 16818 12850 16830
rect 13918 16818 13970 16830
rect 15262 16882 15314 16894
rect 15262 16818 15314 16830
rect 15934 16882 15986 16894
rect 15934 16818 15986 16830
rect 17278 16882 17330 16894
rect 17278 16818 17330 16830
rect 17614 16882 17666 16894
rect 20190 16882 20242 16894
rect 39006 16882 39058 16894
rect 18274 16830 18286 16882
rect 18338 16830 18350 16882
rect 21970 16830 21982 16882
rect 22034 16830 22046 16882
rect 25218 16830 25230 16882
rect 25282 16830 25294 16882
rect 28690 16830 28702 16882
rect 28754 16830 28766 16882
rect 33618 16830 33630 16882
rect 33682 16830 33694 16882
rect 34066 16830 34078 16882
rect 34130 16830 34142 16882
rect 17614 16818 17666 16830
rect 20190 16818 20242 16830
rect 39006 16818 39058 16830
rect 39790 16882 39842 16894
rect 39790 16818 39842 16830
rect 11902 16770 11954 16782
rect 11106 16718 11118 16770
rect 11170 16718 11182 16770
rect 11902 16706 11954 16718
rect 15374 16770 15426 16782
rect 15374 16706 15426 16718
rect 16270 16770 16322 16782
rect 16270 16706 16322 16718
rect 16830 16770 16882 16782
rect 19854 16770 19906 16782
rect 26798 16770 26850 16782
rect 18722 16718 18734 16770
rect 18786 16718 18798 16770
rect 26002 16718 26014 16770
rect 26066 16718 26078 16770
rect 29250 16718 29262 16770
rect 29314 16718 29326 16770
rect 16830 16706 16882 16718
rect 19854 16706 19906 16718
rect 26798 16706 26850 16718
rect 2158 16658 2210 16670
rect 2158 16594 2210 16606
rect 24446 16658 24498 16670
rect 24446 16594 24498 16606
rect 33182 16658 33234 16670
rect 33182 16594 33234 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 10334 16322 10386 16334
rect 10334 16258 10386 16270
rect 12462 16322 12514 16334
rect 12462 16258 12514 16270
rect 12798 16322 12850 16334
rect 12798 16258 12850 16270
rect 13470 16322 13522 16334
rect 13470 16258 13522 16270
rect 18174 16322 18226 16334
rect 18174 16258 18226 16270
rect 34638 16322 34690 16334
rect 34638 16258 34690 16270
rect 36206 16322 36258 16334
rect 36206 16258 36258 16270
rect 12238 16210 12290 16222
rect 12238 16146 12290 16158
rect 13582 16210 13634 16222
rect 13582 16146 13634 16158
rect 14254 16210 14306 16222
rect 20750 16210 20802 16222
rect 31166 16210 31218 16222
rect 35534 16210 35586 16222
rect 19394 16158 19406 16210
rect 19458 16158 19470 16210
rect 26114 16158 26126 16210
rect 26178 16158 26190 16210
rect 32050 16158 32062 16210
rect 32114 16158 32126 16210
rect 14254 16146 14306 16158
rect 20750 16146 20802 16158
rect 31166 16146 31218 16158
rect 35534 16146 35586 16158
rect 36094 16210 36146 16222
rect 36094 16146 36146 16158
rect 14702 16098 14754 16110
rect 21310 16098 21362 16110
rect 28590 16098 28642 16110
rect 2930 16046 2942 16098
rect 2994 16046 3006 16098
rect 6738 16046 6750 16098
rect 6802 16046 6814 16098
rect 7298 16046 7310 16098
rect 7362 16046 7374 16098
rect 15138 16046 15150 16098
rect 15202 16046 15214 16098
rect 19282 16046 19294 16098
rect 19346 16046 19358 16098
rect 21858 16046 21870 16098
rect 21922 16046 21934 16098
rect 25442 16046 25454 16098
rect 25506 16046 25518 16098
rect 14702 16034 14754 16046
rect 21310 16034 21362 16046
rect 28590 16034 28642 16046
rect 29598 16098 29650 16110
rect 29598 16034 29650 16046
rect 31278 16098 31330 16110
rect 31278 16034 31330 16046
rect 31726 16098 31778 16110
rect 34302 16098 34354 16110
rect 32610 16046 32622 16098
rect 32674 16046 32686 16098
rect 32946 16046 32958 16098
rect 33010 16046 33022 16098
rect 33618 16046 33630 16098
rect 33682 16046 33694 16098
rect 38994 16046 39006 16098
rect 39058 16046 39070 16098
rect 31726 16034 31778 16046
rect 34302 16034 34354 16046
rect 12574 15986 12626 15998
rect 2034 15934 2046 15986
rect 2098 15934 2110 15986
rect 12574 15922 12626 15934
rect 19630 15986 19682 15998
rect 19630 15922 19682 15934
rect 25118 15986 25170 15998
rect 25118 15922 25170 15934
rect 27134 15986 27186 15998
rect 27134 15922 27186 15934
rect 27246 15986 27298 15998
rect 27246 15922 27298 15934
rect 28142 15986 28194 15998
rect 31054 15986 31106 15998
rect 29810 15934 29822 15986
rect 29874 15934 29886 15986
rect 30370 15934 30382 15986
rect 30434 15934 30446 15986
rect 28142 15922 28194 15934
rect 31054 15922 31106 15934
rect 33294 15986 33346 15998
rect 33294 15922 33346 15934
rect 33966 15986 34018 15998
rect 33966 15922 34018 15934
rect 34078 15986 34130 15998
rect 34078 15922 34130 15934
rect 34526 15986 34578 15998
rect 40114 15934 40126 15986
rect 40178 15934 40190 15986
rect 34526 15922 34578 15934
rect 10670 15874 10722 15886
rect 26910 15874 26962 15886
rect 9650 15822 9662 15874
rect 9714 15822 9726 15874
rect 17378 15822 17390 15874
rect 17442 15822 17454 15874
rect 24434 15822 24446 15874
rect 24498 15822 24510 15874
rect 10670 15810 10722 15822
rect 26910 15810 26962 15822
rect 27806 15874 27858 15886
rect 27806 15810 27858 15822
rect 29262 15874 29314 15886
rect 29262 15810 29314 15822
rect 32062 15874 32114 15886
rect 32062 15810 32114 15822
rect 32174 15874 32226 15886
rect 32174 15810 32226 15822
rect 32398 15874 32450 15886
rect 32398 15810 32450 15822
rect 33182 15874 33234 15886
rect 33182 15810 33234 15822
rect 33406 15874 33458 15886
rect 33406 15810 33458 15822
rect 35086 15874 35138 15886
rect 35086 15810 35138 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 9662 15538 9714 15550
rect 9662 15474 9714 15486
rect 10110 15538 10162 15550
rect 14142 15538 14194 15550
rect 13570 15486 13582 15538
rect 13634 15486 13646 15538
rect 10110 15474 10162 15486
rect 14142 15474 14194 15486
rect 14366 15538 14418 15550
rect 14366 15474 14418 15486
rect 15598 15538 15650 15550
rect 15598 15474 15650 15486
rect 15822 15538 15874 15550
rect 15822 15474 15874 15486
rect 16830 15538 16882 15550
rect 16830 15474 16882 15486
rect 17502 15538 17554 15550
rect 17502 15474 17554 15486
rect 20078 15538 20130 15550
rect 20078 15474 20130 15486
rect 21758 15538 21810 15550
rect 21758 15474 21810 15486
rect 25790 15538 25842 15550
rect 25790 15474 25842 15486
rect 25902 15538 25954 15550
rect 30270 15538 30322 15550
rect 29474 15486 29486 15538
rect 29538 15486 29550 15538
rect 25902 15474 25954 15486
rect 30270 15474 30322 15486
rect 30718 15538 30770 15550
rect 30718 15474 30770 15486
rect 31614 15538 31666 15550
rect 31614 15474 31666 15486
rect 34638 15538 34690 15550
rect 34638 15474 34690 15486
rect 35534 15538 35586 15550
rect 35534 15474 35586 15486
rect 36094 15538 36146 15550
rect 36094 15474 36146 15486
rect 9550 15426 9602 15438
rect 9550 15362 9602 15374
rect 14478 15426 14530 15438
rect 14478 15362 14530 15374
rect 17614 15426 17666 15438
rect 20862 15426 20914 15438
rect 30494 15426 30546 15438
rect 18498 15374 18510 15426
rect 18562 15374 18574 15426
rect 24098 15374 24110 15426
rect 24162 15374 24174 15426
rect 17614 15362 17666 15374
rect 20862 15362 20914 15374
rect 30494 15362 30546 15374
rect 31950 15426 32002 15438
rect 31950 15362 32002 15374
rect 10670 15314 10722 15326
rect 16270 15314 16322 15326
rect 11106 15262 11118 15314
rect 11170 15262 11182 15314
rect 10670 15250 10722 15262
rect 16270 15250 16322 15262
rect 17278 15314 17330 15326
rect 19182 15314 19234 15326
rect 18722 15262 18734 15314
rect 18786 15262 18798 15314
rect 17278 15250 17330 15262
rect 19182 15250 19234 15262
rect 19406 15314 19458 15326
rect 19406 15250 19458 15262
rect 19630 15314 19682 15326
rect 19630 15250 19682 15262
rect 21758 15314 21810 15326
rect 21758 15250 21810 15262
rect 22094 15314 22146 15326
rect 22094 15250 22146 15262
rect 23326 15314 23378 15326
rect 25678 15314 25730 15326
rect 23762 15262 23774 15314
rect 23826 15262 23838 15314
rect 23326 15250 23378 15262
rect 25678 15250 25730 15262
rect 26350 15314 26402 15326
rect 30942 15314 30994 15326
rect 26674 15262 26686 15314
rect 26738 15262 26750 15314
rect 27234 15262 27246 15314
rect 27298 15262 27310 15314
rect 26350 15250 26402 15262
rect 30942 15250 30994 15262
rect 31054 15314 31106 15326
rect 31054 15250 31106 15262
rect 33294 15314 33346 15326
rect 33294 15250 33346 15262
rect 33630 15314 33682 15326
rect 33630 15250 33682 15262
rect 33854 15314 33906 15326
rect 33854 15250 33906 15262
rect 34078 15314 34130 15326
rect 39006 15314 39058 15326
rect 34402 15262 34414 15314
rect 34466 15262 34478 15314
rect 34078 15250 34130 15262
rect 39006 15250 39058 15262
rect 15374 15202 15426 15214
rect 15374 15138 15426 15150
rect 15710 15202 15762 15214
rect 15710 15138 15762 15150
rect 16718 15202 16770 15214
rect 16718 15138 16770 15150
rect 18062 15202 18114 15214
rect 18062 15138 18114 15150
rect 23214 15202 23266 15214
rect 25230 15202 25282 15214
rect 24434 15150 24446 15202
rect 24498 15150 24510 15202
rect 23214 15138 23266 15150
rect 25230 15138 25282 15150
rect 30830 15202 30882 15214
rect 30830 15138 30882 15150
rect 31502 15202 31554 15214
rect 31502 15138 31554 15150
rect 32510 15202 32562 15214
rect 32510 15138 32562 15150
rect 33406 15202 33458 15214
rect 33406 15138 33458 15150
rect 35086 15202 35138 15214
rect 40350 15202 40402 15214
rect 39778 15150 39790 15202
rect 39842 15150 39854 15202
rect 35086 15138 35138 15150
rect 40350 15138 40402 15150
rect 17950 15090 18002 15102
rect 17950 15026 18002 15038
rect 25342 15090 25394 15102
rect 25342 15026 25394 15038
rect 32062 15090 32114 15102
rect 32062 15026 32114 15038
rect 34750 15090 34802 15102
rect 34750 15026 34802 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 19854 14754 19906 14766
rect 19854 14690 19906 14702
rect 27918 14754 27970 14766
rect 27918 14690 27970 14702
rect 14142 14642 14194 14654
rect 14142 14578 14194 14590
rect 14702 14642 14754 14654
rect 14702 14578 14754 14590
rect 19070 14642 19122 14654
rect 19070 14578 19122 14590
rect 27134 14642 27186 14654
rect 27134 14578 27186 14590
rect 27806 14642 27858 14654
rect 27806 14578 27858 14590
rect 31950 14642 32002 14654
rect 34626 14590 34638 14642
rect 34690 14590 34702 14642
rect 39218 14590 39230 14642
rect 39282 14590 39294 14642
rect 31950 14578 32002 14590
rect 13694 14530 13746 14542
rect 19630 14530 19682 14542
rect 14914 14478 14926 14530
rect 14978 14478 14990 14530
rect 15474 14478 15486 14530
rect 15538 14478 15550 14530
rect 13694 14466 13746 14478
rect 19630 14466 19682 14478
rect 20190 14530 20242 14542
rect 20190 14466 20242 14478
rect 21870 14530 21922 14542
rect 23998 14530 24050 14542
rect 22194 14478 22206 14530
rect 22258 14478 22270 14530
rect 21870 14466 21922 14478
rect 23998 14466 24050 14478
rect 24334 14530 24386 14542
rect 27246 14530 27298 14542
rect 26114 14478 26126 14530
rect 26178 14478 26190 14530
rect 26786 14478 26798 14530
rect 26850 14478 26862 14530
rect 24334 14466 24386 14478
rect 27246 14466 27298 14478
rect 27358 14530 27410 14542
rect 30046 14530 30098 14542
rect 29698 14478 29710 14530
rect 29762 14478 29774 14530
rect 27358 14466 27410 14478
rect 30046 14466 30098 14478
rect 30606 14530 30658 14542
rect 30930 14478 30942 14530
rect 30994 14478 31006 14530
rect 34178 14478 34190 14530
rect 34242 14478 34254 14530
rect 40226 14478 40238 14530
rect 40290 14478 40302 14530
rect 30606 14466 30658 14478
rect 7534 14418 7586 14430
rect 7534 14354 7586 14366
rect 8430 14418 8482 14430
rect 8430 14354 8482 14366
rect 18622 14418 18674 14430
rect 18622 14354 18674 14366
rect 21310 14418 21362 14430
rect 21310 14354 21362 14366
rect 21646 14418 21698 14430
rect 24782 14418 24834 14430
rect 22530 14366 22542 14418
rect 22594 14366 22606 14418
rect 22866 14366 22878 14418
rect 22930 14366 22942 14418
rect 21646 14354 21698 14366
rect 24782 14354 24834 14366
rect 26462 14418 26514 14430
rect 26462 14354 26514 14366
rect 28254 14418 28306 14430
rect 28254 14354 28306 14366
rect 30158 14418 30210 14430
rect 30158 14354 30210 14366
rect 30494 14418 30546 14430
rect 30494 14354 30546 14366
rect 32734 14418 32786 14430
rect 32734 14354 32786 14366
rect 32846 14418 32898 14430
rect 32846 14354 32898 14366
rect 32958 14418 33010 14430
rect 32958 14354 33010 14366
rect 7422 14306 7474 14318
rect 7422 14242 7474 14254
rect 7646 14306 7698 14318
rect 7646 14242 7698 14254
rect 7870 14306 7922 14318
rect 7870 14242 7922 14254
rect 8318 14306 8370 14318
rect 21534 14306 21586 14318
rect 17938 14254 17950 14306
rect 18002 14254 18014 14306
rect 8318 14242 8370 14254
rect 21534 14242 21586 14254
rect 24222 14306 24274 14318
rect 24222 14242 24274 14254
rect 26350 14306 26402 14318
rect 26350 14242 26402 14254
rect 27022 14306 27074 14318
rect 27022 14242 27074 14254
rect 28366 14306 28418 14318
rect 28366 14242 28418 14254
rect 28590 14306 28642 14318
rect 35646 14306 35698 14318
rect 33394 14254 33406 14306
rect 33458 14254 33470 14306
rect 28590 14242 28642 14254
rect 35646 14242 35698 14254
rect 36094 14306 36146 14318
rect 36094 14242 36146 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 16830 13970 16882 13982
rect 21086 13970 21138 13982
rect 26574 13970 26626 13982
rect 19282 13918 19294 13970
rect 19346 13918 19358 13970
rect 24098 13918 24110 13970
rect 24162 13918 24174 13970
rect 16830 13906 16882 13918
rect 21086 13906 21138 13918
rect 26574 13906 26626 13918
rect 33182 13970 33234 13982
rect 33182 13906 33234 13918
rect 38558 13970 38610 13982
rect 38558 13906 38610 13918
rect 5070 13858 5122 13870
rect 16382 13858 16434 13870
rect 8194 13806 8206 13858
rect 8258 13806 8270 13858
rect 13682 13806 13694 13858
rect 13746 13806 13758 13858
rect 5070 13794 5122 13806
rect 16382 13794 16434 13806
rect 17838 13858 17890 13870
rect 20638 13858 20690 13870
rect 19618 13806 19630 13858
rect 19682 13806 19694 13858
rect 17838 13794 17890 13806
rect 20638 13794 20690 13806
rect 22654 13858 22706 13870
rect 22654 13794 22706 13806
rect 27358 13858 27410 13870
rect 27358 13794 27410 13806
rect 28142 13858 28194 13870
rect 32510 13858 32562 13870
rect 30034 13806 30046 13858
rect 30098 13806 30110 13858
rect 30706 13806 30718 13858
rect 30770 13806 30782 13858
rect 28142 13794 28194 13806
rect 32510 13794 32562 13806
rect 33070 13858 33122 13870
rect 33070 13794 33122 13806
rect 33630 13858 33682 13870
rect 33630 13794 33682 13806
rect 37774 13858 37826 13870
rect 37774 13794 37826 13806
rect 5406 13746 5458 13758
rect 21198 13746 21250 13758
rect 8978 13694 8990 13746
rect 9042 13694 9054 13746
rect 15922 13694 15934 13746
rect 15986 13694 15998 13746
rect 19058 13694 19070 13746
rect 19122 13694 19134 13746
rect 20402 13694 20414 13746
rect 20466 13694 20478 13746
rect 5406 13682 5458 13694
rect 21198 13682 21250 13694
rect 21646 13746 21698 13758
rect 21646 13682 21698 13694
rect 22206 13746 22258 13758
rect 26238 13746 26290 13758
rect 27022 13746 27074 13758
rect 25890 13694 25902 13746
rect 25954 13694 25966 13746
rect 26786 13694 26798 13746
rect 26850 13694 26862 13746
rect 22206 13682 22258 13694
rect 26238 13682 26290 13694
rect 27022 13682 27074 13694
rect 27246 13746 27298 13758
rect 27246 13682 27298 13694
rect 27694 13746 27746 13758
rect 27694 13682 27746 13694
rect 28254 13746 28306 13758
rect 31614 13746 31666 13758
rect 28914 13694 28926 13746
rect 28978 13694 28990 13746
rect 30258 13694 30270 13746
rect 30322 13694 30334 13746
rect 31042 13694 31054 13746
rect 31106 13694 31118 13746
rect 28254 13682 28306 13694
rect 31614 13682 31666 13694
rect 32062 13746 32114 13758
rect 32062 13682 32114 13694
rect 32286 13746 32338 13758
rect 32286 13682 32338 13694
rect 33406 13746 33458 13758
rect 34862 13746 34914 13758
rect 34066 13694 34078 13746
rect 34130 13694 34142 13746
rect 35522 13694 35534 13746
rect 35586 13694 35598 13746
rect 38994 13694 39006 13746
rect 39058 13694 39070 13746
rect 33406 13682 33458 13694
rect 34862 13682 34914 13694
rect 9662 13634 9714 13646
rect 6066 13582 6078 13634
rect 6130 13582 6142 13634
rect 9662 13570 9714 13582
rect 21422 13634 21474 13646
rect 21422 13570 21474 13582
rect 23886 13634 23938 13646
rect 27918 13634 27970 13646
rect 32398 13634 32450 13646
rect 25442 13582 25454 13634
rect 25506 13582 25518 13634
rect 27346 13582 27358 13634
rect 27410 13582 27422 13634
rect 31154 13582 31166 13634
rect 31218 13582 31230 13634
rect 34514 13582 34526 13634
rect 34578 13582 34590 13634
rect 40002 13582 40014 13634
rect 40066 13582 40078 13634
rect 23886 13570 23938 13582
rect 27918 13570 27970 13582
rect 32398 13570 32450 13582
rect 21086 13522 21138 13534
rect 21086 13458 21138 13470
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 7198 13186 7250 13198
rect 7198 13122 7250 13134
rect 7310 13186 7362 13198
rect 7310 13122 7362 13134
rect 7534 13186 7586 13198
rect 7534 13122 7586 13134
rect 18846 13186 18898 13198
rect 26910 13186 26962 13198
rect 26002 13134 26014 13186
rect 26066 13134 26078 13186
rect 18846 13122 18898 13134
rect 26910 13122 26962 13134
rect 30158 13186 30210 13198
rect 32510 13186 32562 13198
rect 31266 13134 31278 13186
rect 31330 13183 31342 13186
rect 31826 13183 31838 13186
rect 31330 13137 31838 13183
rect 31330 13134 31342 13137
rect 31826 13134 31838 13137
rect 31890 13134 31902 13186
rect 30158 13122 30210 13134
rect 32510 13122 32562 13134
rect 32734 13186 32786 13198
rect 32734 13122 32786 13134
rect 37774 13186 37826 13198
rect 37774 13122 37826 13134
rect 5630 13074 5682 13086
rect 12014 13074 12066 13086
rect 2930 13022 2942 13074
rect 2994 13022 3006 13074
rect 5058 13022 5070 13074
rect 5122 13022 5134 13074
rect 6514 13022 6526 13074
rect 6578 13022 6590 13074
rect 10882 13022 10894 13074
rect 10946 13022 10958 13074
rect 5630 13010 5682 13022
rect 12014 13010 12066 13022
rect 12462 13074 12514 13086
rect 12462 13010 12514 13022
rect 12910 13074 12962 13086
rect 12910 13010 12962 13022
rect 13694 13074 13746 13086
rect 21646 13074 21698 13086
rect 27134 13074 27186 13086
rect 15250 13022 15262 13074
rect 15314 13022 15326 13074
rect 18498 13022 18510 13074
rect 18562 13022 18574 13074
rect 20402 13022 20414 13074
rect 20466 13022 20478 13074
rect 22866 13022 22878 13074
rect 22930 13022 22942 13074
rect 13694 13010 13746 13022
rect 21646 13010 21698 13022
rect 27134 13010 27186 13022
rect 29262 13074 29314 13086
rect 29262 13010 29314 13022
rect 31502 13074 31554 13086
rect 31502 13010 31554 13022
rect 31950 13074 32002 13086
rect 31950 13010 32002 13022
rect 34190 13074 34242 13086
rect 34190 13010 34242 13022
rect 37326 13074 37378 13086
rect 37326 13010 37378 13022
rect 37662 13074 37714 13086
rect 37662 13010 37714 13022
rect 38670 13074 38722 13086
rect 38670 13010 38722 13022
rect 19070 12962 19122 12974
rect 2258 12910 2270 12962
rect 2322 12910 2334 12962
rect 6066 12910 6078 12962
rect 6130 12910 6142 12962
rect 7970 12910 7982 12962
rect 8034 12910 8046 12962
rect 19070 12898 19122 12910
rect 19406 12962 19458 12974
rect 19406 12898 19458 12910
rect 19742 12962 19794 12974
rect 26686 12962 26738 12974
rect 28030 12962 28082 12974
rect 20626 12910 20638 12962
rect 20690 12910 20702 12962
rect 22082 12910 22094 12962
rect 22146 12910 22158 12962
rect 23650 12910 23662 12962
rect 23714 12910 23726 12962
rect 24770 12910 24782 12962
rect 24834 12910 24846 12962
rect 25218 12910 25230 12962
rect 25282 12910 25294 12962
rect 27794 12910 27806 12962
rect 27858 12910 27870 12962
rect 19742 12898 19794 12910
rect 26686 12898 26738 12910
rect 28030 12898 28082 12910
rect 28366 12962 28418 12974
rect 28366 12898 28418 12910
rect 29150 12962 29202 12974
rect 29150 12898 29202 12910
rect 29822 12962 29874 12974
rect 29822 12898 29874 12910
rect 30046 12962 30098 12974
rect 33182 12962 33234 12974
rect 33058 12910 33070 12962
rect 33122 12910 33134 12962
rect 30046 12898 30098 12910
rect 33182 12898 33234 12910
rect 33406 12962 33458 12974
rect 33406 12898 33458 12910
rect 34078 12962 34130 12974
rect 34078 12898 34130 12910
rect 34750 12962 34802 12974
rect 34750 12898 34802 12910
rect 35310 12962 35362 12974
rect 35310 12898 35362 12910
rect 35758 12962 35810 12974
rect 35758 12898 35810 12910
rect 35982 12962 36034 12974
rect 35982 12898 36034 12910
rect 7646 12850 7698 12862
rect 11230 12850 11282 12862
rect 18286 12850 18338 12862
rect 8754 12798 8766 12850
rect 8818 12798 8830 12850
rect 14354 12798 14366 12850
rect 14418 12798 14430 12850
rect 7646 12786 7698 12798
rect 11230 12786 11282 12798
rect 18286 12786 18338 12798
rect 18510 12850 18562 12862
rect 27582 12850 27634 12862
rect 20402 12798 20414 12850
rect 20466 12798 20478 12850
rect 18510 12786 18562 12798
rect 27582 12786 27634 12798
rect 30830 12850 30882 12862
rect 30830 12786 30882 12798
rect 34974 12850 35026 12862
rect 34974 12786 35026 12798
rect 35646 12850 35698 12862
rect 35646 12786 35698 12798
rect 36318 12850 36370 12862
rect 36318 12786 36370 12798
rect 39454 12850 39506 12862
rect 39454 12786 39506 12798
rect 39678 12850 39730 12862
rect 39678 12786 39730 12798
rect 40238 12850 40290 12862
rect 40238 12786 40290 12798
rect 11342 12738 11394 12750
rect 11342 12674 11394 12686
rect 11454 12738 11506 12750
rect 11454 12674 11506 12686
rect 11902 12738 11954 12750
rect 11902 12674 11954 12686
rect 19630 12738 19682 12750
rect 19630 12674 19682 12686
rect 28142 12738 28194 12750
rect 28142 12674 28194 12686
rect 28254 12738 28306 12750
rect 28254 12674 28306 12686
rect 29374 12738 29426 12750
rect 29374 12674 29426 12686
rect 30158 12738 30210 12750
rect 30158 12674 30210 12686
rect 30942 12738 30994 12750
rect 30942 12674 30994 12686
rect 31166 12738 31218 12750
rect 31166 12674 31218 12686
rect 33294 12738 33346 12750
rect 33294 12674 33346 12686
rect 34302 12738 34354 12750
rect 34302 12674 34354 12686
rect 35086 12738 35138 12750
rect 35086 12674 35138 12686
rect 35422 12738 35474 12750
rect 35422 12674 35474 12686
rect 36206 12738 36258 12750
rect 36206 12674 36258 12686
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 4846 12402 4898 12414
rect 4846 12338 4898 12350
rect 18286 12402 18338 12414
rect 18286 12338 18338 12350
rect 20974 12402 21026 12414
rect 20974 12338 21026 12350
rect 27582 12402 27634 12414
rect 32398 12402 32450 12414
rect 30706 12350 30718 12402
rect 30770 12350 30782 12402
rect 27582 12338 27634 12350
rect 32398 12338 32450 12350
rect 34526 12402 34578 12414
rect 34526 12338 34578 12350
rect 8542 12290 8594 12302
rect 18846 12290 18898 12302
rect 14690 12238 14702 12290
rect 14754 12238 14766 12290
rect 8542 12226 8594 12238
rect 18846 12226 18898 12238
rect 19294 12290 19346 12302
rect 25790 12290 25842 12302
rect 34974 12290 35026 12302
rect 21970 12238 21982 12290
rect 22034 12238 22046 12290
rect 22978 12238 22990 12290
rect 23042 12238 23054 12290
rect 28914 12238 28926 12290
rect 28978 12238 28990 12290
rect 30594 12238 30606 12290
rect 30658 12238 30670 12290
rect 31266 12238 31278 12290
rect 31330 12238 31342 12290
rect 33730 12238 33742 12290
rect 33794 12238 33806 12290
rect 19294 12226 19346 12238
rect 25790 12226 25842 12238
rect 34974 12226 35026 12238
rect 17950 12178 18002 12190
rect 30494 12178 30546 12190
rect 34750 12178 34802 12190
rect 5170 12126 5182 12178
rect 5234 12126 5246 12178
rect 13458 12126 13470 12178
rect 13522 12126 13534 12178
rect 13906 12126 13918 12178
rect 13970 12126 13982 12178
rect 19954 12126 19966 12178
rect 20018 12126 20030 12178
rect 20850 12126 20862 12178
rect 20914 12126 20926 12178
rect 22194 12126 22206 12178
rect 22258 12126 22270 12178
rect 23090 12126 23102 12178
rect 23154 12126 23166 12178
rect 25218 12126 25230 12178
rect 25282 12126 25294 12178
rect 28466 12126 28478 12178
rect 28530 12126 28542 12178
rect 29474 12126 29486 12178
rect 29538 12126 29550 12178
rect 30034 12126 30046 12178
rect 30098 12126 30110 12178
rect 33058 12126 33070 12178
rect 33122 12126 33134 12178
rect 33618 12126 33630 12178
rect 33682 12126 33694 12178
rect 17950 12114 18002 12126
rect 30494 12114 30546 12126
rect 34750 12114 34802 12126
rect 18398 12066 18450 12078
rect 27022 12066 27074 12078
rect 34638 12066 34690 12078
rect 5954 12014 5966 12066
rect 6018 12014 6030 12066
rect 8082 12014 8094 12066
rect 8146 12014 8158 12066
rect 10658 12014 10670 12066
rect 10722 12014 10734 12066
rect 12786 12014 12798 12066
rect 12850 12014 12862 12066
rect 16818 12014 16830 12066
rect 16882 12014 16894 12066
rect 20738 12014 20750 12066
rect 20802 12014 20814 12066
rect 22754 12014 22766 12066
rect 22818 12014 22830 12066
rect 28802 12014 28814 12066
rect 28866 12014 28878 12066
rect 34066 12014 34078 12066
rect 34130 12014 34142 12066
rect 18398 12002 18450 12014
rect 27022 12002 27074 12014
rect 34638 12002 34690 12014
rect 35534 12066 35586 12078
rect 35534 12002 35586 12014
rect 35982 12066 36034 12078
rect 35982 12002 36034 12014
rect 17726 11954 17778 11966
rect 17378 11902 17390 11954
rect 17442 11902 17454 11954
rect 17726 11890 17778 11902
rect 18734 11954 18786 11966
rect 18734 11890 18786 11902
rect 19854 11954 19906 11966
rect 19854 11890 19906 11902
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 6862 11618 6914 11630
rect 6862 11554 6914 11566
rect 27246 11618 27298 11630
rect 27246 11554 27298 11566
rect 27806 11618 27858 11630
rect 27806 11554 27858 11566
rect 28254 11618 28306 11630
rect 28254 11554 28306 11566
rect 6974 11506 7026 11518
rect 27358 11506 27410 11518
rect 12898 11454 12910 11506
rect 12962 11454 12974 11506
rect 20514 11454 20526 11506
rect 20578 11454 20590 11506
rect 22642 11454 22654 11506
rect 22706 11454 22718 11506
rect 25330 11454 25342 11506
rect 25394 11454 25406 11506
rect 6974 11442 7026 11454
rect 27358 11442 27410 11454
rect 27694 11506 27746 11518
rect 27694 11442 27746 11454
rect 29710 11506 29762 11518
rect 29710 11442 29762 11454
rect 13582 11394 13634 11406
rect 14926 11394 14978 11406
rect 27918 11394 27970 11406
rect 9426 11342 9438 11394
rect 9490 11342 9502 11394
rect 9986 11342 9998 11394
rect 10050 11342 10062 11394
rect 13906 11342 13918 11394
rect 13970 11342 13982 11394
rect 15586 11342 15598 11394
rect 15650 11342 15662 11394
rect 20402 11342 20414 11394
rect 20466 11342 20478 11394
rect 22866 11342 22878 11394
rect 22930 11342 22942 11394
rect 23762 11342 23774 11394
rect 23826 11342 23838 11394
rect 25442 11342 25454 11394
rect 25506 11342 25518 11394
rect 13582 11330 13634 11342
rect 14926 11330 14978 11342
rect 27918 11330 27970 11342
rect 28478 11394 28530 11406
rect 28478 11330 28530 11342
rect 29598 11394 29650 11406
rect 29598 11330 29650 11342
rect 29934 11394 29986 11406
rect 29934 11330 29986 11342
rect 30046 11394 30098 11406
rect 31166 11394 31218 11406
rect 34190 11394 34242 11406
rect 30482 11342 30494 11394
rect 30546 11342 30558 11394
rect 32050 11342 32062 11394
rect 32114 11342 32126 11394
rect 32834 11342 32846 11394
rect 32898 11342 32910 11394
rect 33394 11342 33406 11394
rect 33458 11342 33470 11394
rect 30046 11330 30098 11342
rect 31166 11330 31218 11342
rect 34190 11330 34242 11342
rect 34526 11394 34578 11406
rect 34526 11330 34578 11342
rect 34750 11394 34802 11406
rect 35870 11394 35922 11406
rect 35634 11342 35646 11394
rect 35698 11342 35710 11394
rect 34750 11330 34802 11342
rect 35870 11330 35922 11342
rect 36206 11394 36258 11406
rect 36206 11330 36258 11342
rect 13470 11282 13522 11294
rect 10770 11230 10782 11282
rect 10834 11230 10846 11282
rect 13470 11218 13522 11230
rect 19406 11282 19458 11294
rect 19406 11218 19458 11230
rect 19742 11282 19794 11294
rect 25118 11282 25170 11294
rect 21858 11230 21870 11282
rect 21922 11230 21934 11282
rect 24434 11230 24446 11282
rect 24498 11230 24510 11282
rect 19742 11218 19794 11230
rect 25118 11218 25170 11230
rect 30942 11282 30994 11294
rect 30942 11218 30994 11230
rect 31054 11282 31106 11294
rect 31054 11218 31106 11230
rect 31278 11282 31330 11294
rect 35086 11282 35138 11294
rect 31714 11230 31726 11282
rect 31778 11230 31790 11282
rect 32722 11230 32734 11282
rect 32786 11230 32798 11282
rect 31278 11218 31330 11230
rect 35086 11218 35138 11230
rect 36094 11282 36146 11294
rect 36094 11218 36146 11230
rect 37214 11282 37266 11294
rect 37214 11218 37266 11230
rect 9662 11170 9714 11182
rect 18622 11170 18674 11182
rect 18050 11118 18062 11170
rect 18114 11118 18126 11170
rect 9662 11106 9714 11118
rect 18622 11106 18674 11118
rect 19070 11170 19122 11182
rect 19070 11106 19122 11118
rect 29262 11170 29314 11182
rect 29262 11106 29314 11118
rect 33966 11170 34018 11182
rect 33966 11106 34018 11118
rect 34302 11170 34354 11182
rect 34302 11106 34354 11118
rect 35198 11170 35250 11182
rect 35198 11106 35250 11118
rect 35310 11170 35362 11182
rect 35310 11106 35362 11118
rect 37774 11170 37826 11182
rect 37774 11106 37826 11118
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 12798 10834 12850 10846
rect 30046 10834 30098 10846
rect 16706 10782 16718 10834
rect 16770 10782 16782 10834
rect 12798 10770 12850 10782
rect 30046 10770 30098 10782
rect 30382 10834 30434 10846
rect 30382 10770 30434 10782
rect 31278 10834 31330 10846
rect 31278 10770 31330 10782
rect 31502 10834 31554 10846
rect 38334 10834 38386 10846
rect 37762 10782 37774 10834
rect 37826 10782 37838 10834
rect 31502 10770 31554 10782
rect 38334 10770 38386 10782
rect 13134 10722 13186 10734
rect 10322 10670 10334 10722
rect 10386 10670 10398 10722
rect 13134 10658 13186 10670
rect 17502 10722 17554 10734
rect 17502 10658 17554 10670
rect 17838 10722 17890 10734
rect 17838 10658 17890 10670
rect 20974 10722 21026 10734
rect 27022 10722 27074 10734
rect 25330 10670 25342 10722
rect 25394 10670 25406 10722
rect 20974 10658 21026 10670
rect 27022 10658 27074 10670
rect 27134 10722 27186 10734
rect 30494 10722 30546 10734
rect 28130 10670 28142 10722
rect 28194 10670 28206 10722
rect 28802 10670 28814 10722
rect 28866 10670 28878 10722
rect 27134 10658 27186 10670
rect 30494 10658 30546 10670
rect 31614 10722 31666 10734
rect 31614 10658 31666 10670
rect 32062 10722 32114 10734
rect 32062 10658 32114 10670
rect 33070 10722 33122 10734
rect 33070 10658 33122 10670
rect 38670 10722 38722 10734
rect 38670 10658 38722 10670
rect 39118 10722 39170 10734
rect 39118 10658 39170 10670
rect 32286 10610 32338 10622
rect 9650 10558 9662 10610
rect 9714 10558 9726 10610
rect 13682 10558 13694 10610
rect 13746 10558 13758 10610
rect 18162 10558 18174 10610
rect 18226 10558 18238 10610
rect 18722 10558 18734 10610
rect 18786 10558 18798 10610
rect 25218 10558 25230 10610
rect 25282 10558 25294 10610
rect 27346 10558 27358 10610
rect 27410 10558 27422 10610
rect 28018 10558 28030 10610
rect 28082 10558 28094 10610
rect 28914 10558 28926 10610
rect 28978 10558 28990 10610
rect 29922 10558 29934 10610
rect 29986 10558 29998 10610
rect 32286 10546 32338 10558
rect 32510 10610 32562 10622
rect 33966 10610 34018 10622
rect 33730 10558 33742 10610
rect 33794 10558 33806 10610
rect 32510 10546 32562 10558
rect 33966 10546 34018 10558
rect 34862 10610 34914 10622
rect 38558 10610 38610 10622
rect 35298 10558 35310 10610
rect 35362 10558 35374 10610
rect 34862 10546 34914 10558
rect 38558 10546 38610 10558
rect 22206 10498 22258 10510
rect 30942 10498 30994 10510
rect 12450 10446 12462 10498
rect 12514 10446 12526 10498
rect 14466 10446 14478 10498
rect 14530 10446 14542 10498
rect 25890 10446 25902 10498
rect 25954 10446 25966 10498
rect 22206 10434 22258 10446
rect 30942 10434 30994 10446
rect 32398 10498 32450 10510
rect 32398 10434 32450 10446
rect 26562 10334 26574 10386
rect 26626 10334 26638 10386
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 11118 10050 11170 10062
rect 10770 9998 10782 10050
rect 10834 9998 10846 10050
rect 11118 9986 11170 9998
rect 14814 10050 14866 10062
rect 14814 9986 14866 9998
rect 19742 10050 19794 10062
rect 19742 9986 19794 9998
rect 29150 10050 29202 10062
rect 29150 9986 29202 9998
rect 29710 10050 29762 10062
rect 29710 9986 29762 9998
rect 29934 10050 29986 10062
rect 29934 9986 29986 9998
rect 34638 10050 34690 10062
rect 34638 9986 34690 9998
rect 11342 9938 11394 9950
rect 11342 9874 11394 9886
rect 12574 9938 12626 9950
rect 12574 9874 12626 9886
rect 13022 9938 13074 9950
rect 13022 9874 13074 9886
rect 13694 9938 13746 9950
rect 13694 9874 13746 9886
rect 13918 9938 13970 9950
rect 13918 9874 13970 9886
rect 15374 9938 15426 9950
rect 15374 9874 15426 9886
rect 19294 9938 19346 9950
rect 19294 9874 19346 9886
rect 19630 9938 19682 9950
rect 20514 9886 20526 9938
rect 20578 9886 20590 9938
rect 21634 9886 21646 9938
rect 21698 9886 21710 9938
rect 22306 9886 22318 9938
rect 22370 9886 22382 9938
rect 19630 9874 19682 9886
rect 24334 9826 24386 9838
rect 20738 9774 20750 9826
rect 20802 9774 20814 9826
rect 21298 9774 21310 9826
rect 21362 9774 21374 9826
rect 22418 9774 22430 9826
rect 22482 9774 22494 9826
rect 24334 9762 24386 9774
rect 24782 9826 24834 9838
rect 24782 9762 24834 9774
rect 25006 9826 25058 9838
rect 30382 9826 30434 9838
rect 26562 9774 26574 9826
rect 26626 9774 26638 9826
rect 25006 9762 25058 9774
rect 30382 9762 30434 9774
rect 30606 9826 30658 9838
rect 32834 9774 32846 9826
rect 32898 9774 32910 9826
rect 30606 9762 30658 9774
rect 14478 9714 14530 9726
rect 20514 9662 20526 9714
rect 20578 9662 20590 9714
rect 23090 9673 23102 9725
rect 23154 9673 23166 9725
rect 28478 9714 28530 9726
rect 26002 9662 26014 9714
rect 26066 9662 26078 9714
rect 27682 9662 27694 9714
rect 27746 9662 27758 9714
rect 14478 9650 14530 9662
rect 28478 9650 28530 9662
rect 28590 9714 28642 9726
rect 28590 9650 28642 9662
rect 29374 9714 29426 9726
rect 34638 9714 34690 9726
rect 32274 9662 32286 9714
rect 32338 9662 32350 9714
rect 33954 9662 33966 9714
rect 34018 9662 34030 9714
rect 29374 9650 29426 9662
rect 34638 9650 34690 9662
rect 34750 9658 34802 9670
rect 14030 9602 14082 9614
rect 14030 9538 14082 9550
rect 14702 9602 14754 9614
rect 14702 9538 14754 9550
rect 24894 9602 24946 9614
rect 24894 9538 24946 9550
rect 25230 9602 25282 9614
rect 28254 9602 28306 9614
rect 27794 9550 27806 9602
rect 27858 9550 27870 9602
rect 25230 9538 25282 9550
rect 28254 9538 28306 9550
rect 30046 9602 30098 9614
rect 30046 9538 30098 9550
rect 30494 9602 30546 9614
rect 30494 9538 30546 9550
rect 30830 9602 30882 9614
rect 30830 9538 30882 9550
rect 31390 9602 31442 9614
rect 33842 9550 33854 9602
rect 33906 9550 33918 9602
rect 34750 9594 34802 9606
rect 35310 9602 35362 9614
rect 31390 9538 31442 9550
rect 35310 9538 35362 9550
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 21870 9266 21922 9278
rect 24782 9266 24834 9278
rect 21298 9214 21310 9266
rect 21362 9214 21374 9266
rect 23202 9214 23214 9266
rect 23266 9214 23278 9266
rect 21870 9202 21922 9214
rect 24782 9202 24834 9214
rect 26798 9266 26850 9278
rect 26798 9202 26850 9214
rect 27358 9266 27410 9278
rect 27358 9202 27410 9214
rect 27582 9266 27634 9278
rect 31950 9266 32002 9278
rect 30370 9214 30382 9266
rect 30434 9214 30446 9266
rect 27582 9202 27634 9214
rect 31950 9202 32002 9214
rect 32174 9266 32226 9278
rect 32174 9202 32226 9214
rect 33406 9266 33458 9278
rect 33406 9202 33458 9214
rect 34078 9266 34130 9278
rect 34078 9202 34130 9214
rect 34638 9266 34690 9278
rect 34638 9202 34690 9214
rect 35086 9266 35138 9278
rect 35086 9202 35138 9214
rect 27022 9154 27074 9166
rect 26002 9102 26014 9154
rect 26066 9102 26078 9154
rect 26450 9102 26462 9154
rect 26514 9102 26526 9154
rect 27022 9090 27074 9102
rect 27134 9154 27186 9166
rect 27134 9090 27186 9102
rect 27694 9154 27746 9166
rect 31502 9154 31554 9166
rect 28578 9102 28590 9154
rect 28642 9102 28654 9154
rect 30258 9102 30270 9154
rect 30322 9102 30334 9154
rect 27694 9090 27746 9102
rect 31502 9090 31554 9102
rect 33854 9154 33906 9166
rect 33854 9090 33906 9102
rect 34190 9154 34242 9166
rect 34190 9090 34242 9102
rect 18174 9042 18226 9054
rect 25678 9042 25730 9054
rect 31614 9042 31666 9054
rect 18834 8990 18846 9042
rect 18898 8990 18910 9042
rect 22418 8990 22430 9042
rect 22482 8990 22494 9042
rect 22642 8990 22654 9042
rect 22706 8990 22718 9042
rect 22866 8990 22878 9042
rect 22930 8990 22942 9042
rect 29138 8990 29150 9042
rect 29202 8990 29214 9042
rect 18174 8978 18226 8990
rect 25678 8978 25730 8990
rect 31614 8978 31666 8990
rect 32062 9042 32114 9054
rect 32062 8978 32114 8990
rect 32622 9042 32674 9054
rect 32622 8978 32674 8990
rect 33070 9042 33122 9054
rect 33070 8978 33122 8990
rect 33406 9042 33458 9054
rect 33406 8978 33458 8990
rect 33742 9042 33794 9054
rect 33742 8978 33794 8990
rect 30942 8930 30994 8942
rect 30942 8866 30994 8878
rect 25342 8818 25394 8830
rect 25342 8754 25394 8766
rect 31502 8818 31554 8830
rect 31502 8754 31554 8766
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 21310 8482 21362 8494
rect 21310 8418 21362 8430
rect 25678 8482 25730 8494
rect 25678 8418 25730 8430
rect 21422 8370 21474 8382
rect 20626 8318 20638 8370
rect 20690 8318 20702 8370
rect 21422 8306 21474 8318
rect 30158 8370 30210 8382
rect 30158 8306 30210 8318
rect 30606 8370 30658 8382
rect 30606 8306 30658 8318
rect 31166 8370 31218 8382
rect 31166 8306 31218 8318
rect 31726 8370 31778 8382
rect 31726 8306 31778 8318
rect 32174 8370 32226 8382
rect 32174 8306 32226 8318
rect 36318 8370 36370 8382
rect 36318 8306 36370 8318
rect 22206 8258 22258 8270
rect 28254 8258 28306 8270
rect 20402 8206 20414 8258
rect 20466 8206 20478 8258
rect 22642 8206 22654 8258
rect 22706 8206 22718 8258
rect 26338 8206 26350 8258
rect 26402 8206 26414 8258
rect 22206 8194 22258 8206
rect 28254 8194 28306 8206
rect 29150 8258 29202 8270
rect 29150 8194 29202 8206
rect 29374 8258 29426 8270
rect 32622 8258 32674 8270
rect 29698 8206 29710 8258
rect 29762 8206 29774 8258
rect 33170 8206 33182 8258
rect 33234 8206 33246 8258
rect 29374 8194 29426 8206
rect 32622 8194 32674 8206
rect 19406 8146 19458 8158
rect 19406 8082 19458 8094
rect 19742 8146 19794 8158
rect 19742 8082 19794 8094
rect 26014 8146 26066 8158
rect 28030 8146 28082 8158
rect 27458 8094 27470 8146
rect 27522 8094 27534 8146
rect 26014 8082 26066 8094
rect 28030 8082 28082 8094
rect 28478 8146 28530 8158
rect 28478 8082 28530 8094
rect 28590 8146 28642 8158
rect 28590 8082 28642 8094
rect 19070 8034 19122 8046
rect 25902 8034 25954 8046
rect 25106 7982 25118 8034
rect 25170 7982 25182 8034
rect 19070 7970 19122 7982
rect 25902 7970 25954 7982
rect 27918 8034 27970 8046
rect 27918 7970 27970 7982
rect 29262 8034 29314 8046
rect 35746 7982 35758 8034
rect 35810 7982 35822 8034
rect 29262 7970 29314 7982
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 22318 7698 22370 7710
rect 21298 7646 21310 7698
rect 21362 7646 21374 7698
rect 22318 7634 22370 7646
rect 26238 7698 26290 7710
rect 26238 7634 26290 7646
rect 26910 7698 26962 7710
rect 26910 7634 26962 7646
rect 27470 7698 27522 7710
rect 27470 7634 27522 7646
rect 27918 7698 27970 7710
rect 27918 7634 27970 7646
rect 33182 7698 33234 7710
rect 33182 7634 33234 7646
rect 35758 7698 35810 7710
rect 35758 7634 35810 7646
rect 23438 7586 23490 7598
rect 23438 7522 23490 7534
rect 23774 7586 23826 7598
rect 23774 7522 23826 7534
rect 28702 7586 28754 7598
rect 28702 7522 28754 7534
rect 31838 7586 31890 7598
rect 31838 7522 31890 7534
rect 31950 7586 32002 7598
rect 31950 7522 32002 7534
rect 32398 7586 32450 7598
rect 32398 7522 32450 7534
rect 35422 7586 35474 7598
rect 35422 7522 35474 7534
rect 35870 7586 35922 7598
rect 35870 7522 35922 7534
rect 18174 7474 18226 7486
rect 31390 7474 31442 7486
rect 18834 7422 18846 7474
rect 18898 7422 18910 7474
rect 30930 7422 30942 7474
rect 30994 7422 31006 7474
rect 18174 7410 18226 7422
rect 31390 7410 31442 7422
rect 25790 7362 25842 7374
rect 25790 7298 25842 7310
rect 25554 7198 25566 7250
rect 25618 7247 25630 7250
rect 26450 7247 26462 7250
rect 25618 7201 26462 7247
rect 25618 7198 25630 7201
rect 26450 7198 26462 7201
rect 26514 7198 26526 7250
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 21310 6914 21362 6926
rect 21310 6850 21362 6862
rect 27470 6914 27522 6926
rect 27470 6850 27522 6862
rect 21422 6802 21474 6814
rect 21422 6738 21474 6750
rect 31838 6802 31890 6814
rect 31838 6738 31890 6750
rect 21982 6690 22034 6702
rect 21982 6626 22034 6638
rect 23774 6690 23826 6702
rect 28366 6690 28418 6702
rect 24434 6638 24446 6690
rect 24498 6638 24510 6690
rect 23774 6626 23826 6638
rect 28366 6626 28418 6638
rect 22430 6466 22482 6478
rect 27918 6466 27970 6478
rect 26786 6414 26798 6466
rect 26850 6414 26862 6466
rect 22430 6402 22482 6414
rect 27918 6402 27970 6414
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 17490 4286 17502 4338
rect 17554 4286 17566 4338
rect 26350 4226 26402 4238
rect 17826 4174 17838 4226
rect 17890 4174 17902 4226
rect 26350 4162 26402 4174
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 18834 3614 18846 3666
rect 18898 3614 18910 3666
rect 22194 3614 22206 3666
rect 22258 3614 22270 3666
rect 25666 3614 25678 3666
rect 25730 3614 25742 3666
rect 26898 3614 26910 3666
rect 26962 3614 26974 3666
rect 23102 3554 23154 3566
rect 26126 3554 26178 3566
rect 23538 3502 23550 3554
rect 23602 3502 23614 3554
rect 23102 3490 23154 3502
rect 26126 3490 26178 3502
rect 26462 3554 26514 3566
rect 26462 3490 26514 3502
rect 18398 3442 18450 3454
rect 18398 3378 18450 3390
rect 21758 3442 21810 3454
rect 21758 3378 21810 3390
rect 23326 3442 23378 3454
rect 23326 3378 23378 3390
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 8766 38558 8818 38610
rect 9774 38558 9826 38610
rect 12126 38558 12178 38610
rect 13134 38558 13186 38610
rect 15934 38558 15986 38610
rect 16718 38558 16770 38610
rect 25566 38558 25618 38610
rect 26350 38558 26402 38610
rect 27022 38558 27074 38610
rect 28478 38558 28530 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 13134 38222 13186 38274
rect 15486 38222 15538 38274
rect 18174 38222 18226 38274
rect 20190 38222 20242 38274
rect 9774 38110 9826 38162
rect 12686 38110 12738 38162
rect 18734 38110 18786 38162
rect 21310 38110 21362 38162
rect 22878 38110 22930 38162
rect 24782 38110 24834 38162
rect 26350 38110 26402 38162
rect 28814 38110 28866 38162
rect 30382 38110 30434 38162
rect 32734 38110 32786 38162
rect 34414 38110 34466 38162
rect 11006 37998 11058 38050
rect 11678 37998 11730 38050
rect 17502 37998 17554 38050
rect 22094 37998 22146 38050
rect 23438 37998 23490 38050
rect 25566 37998 25618 38050
rect 27246 37998 27298 38050
rect 28478 37998 28530 38050
rect 33742 37998 33794 38050
rect 35422 37998 35474 38050
rect 9326 37774 9378 37826
rect 11454 37774 11506 37826
rect 12014 37774 12066 37826
rect 13918 37774 13970 37826
rect 14814 37774 14866 37826
rect 15262 37774 15314 37826
rect 16270 37774 16322 37826
rect 17166 37774 17218 37826
rect 19182 37774 19234 37826
rect 19406 37774 19458 37826
rect 23998 37774 24050 37826
rect 27806 37774 27858 37826
rect 29710 37774 29762 37826
rect 29934 37774 29986 37826
rect 31278 37774 31330 37826
rect 31614 37774 31666 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 9102 37438 9154 37490
rect 9662 37438 9714 37490
rect 14590 37438 14642 37490
rect 15934 37438 15986 37490
rect 17390 37438 17442 37490
rect 18958 37438 19010 37490
rect 22654 37438 22706 37490
rect 23214 37438 23266 37490
rect 23998 37438 24050 37490
rect 28926 37438 28978 37490
rect 29598 37438 29650 37490
rect 32398 37438 32450 37490
rect 34974 37438 35026 37490
rect 19294 37326 19346 37378
rect 24334 37326 24386 37378
rect 25230 37326 25282 37378
rect 25342 37326 25394 37378
rect 31390 37326 31442 37378
rect 11678 37214 11730 37266
rect 12126 37214 12178 37266
rect 16718 37214 16770 37266
rect 18062 37214 18114 37266
rect 19518 37214 19570 37266
rect 20190 37214 20242 37266
rect 24670 37214 24722 37266
rect 25566 37214 25618 37266
rect 25902 37214 25954 37266
rect 26574 37214 26626 37266
rect 29822 37214 29874 37266
rect 30270 37214 30322 37266
rect 31166 37214 31218 37266
rect 31502 37214 31554 37266
rect 33630 37214 33682 37266
rect 10110 37102 10162 37154
rect 10782 37102 10834 37154
rect 11230 37102 11282 37154
rect 15486 37102 15538 37154
rect 16382 37102 16434 37154
rect 18622 37102 18674 37154
rect 23438 37102 23490 37154
rect 30830 37102 30882 37154
rect 31950 37102 32002 37154
rect 33294 37102 33346 37154
rect 34078 37102 34130 37154
rect 34526 37102 34578 37154
rect 15150 36990 15202 37042
rect 30942 36990 30994 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 12574 36654 12626 36706
rect 14926 36654 14978 36706
rect 22878 36654 22930 36706
rect 27246 36654 27298 36706
rect 32734 36654 32786 36706
rect 36542 36654 36594 36706
rect 12910 36542 12962 36594
rect 16158 36542 16210 36594
rect 21422 36542 21474 36594
rect 27582 36542 27634 36594
rect 9102 36430 9154 36482
rect 9550 36430 9602 36482
rect 15374 36430 15426 36482
rect 16494 36430 16546 36482
rect 17054 36430 17106 36482
rect 21982 36430 22034 36482
rect 23550 36430 23602 36482
rect 24222 36430 24274 36482
rect 28030 36430 28082 36482
rect 28254 36430 28306 36482
rect 29038 36430 29090 36482
rect 29710 36430 29762 36482
rect 32846 36430 32898 36482
rect 33406 36430 33458 36482
rect 13470 36318 13522 36370
rect 13806 36318 13858 36370
rect 14590 36318 14642 36370
rect 15710 36318 15762 36370
rect 20526 36318 20578 36370
rect 22990 36318 23042 36370
rect 27470 36318 27522 36370
rect 27694 36318 27746 36370
rect 28478 36318 28530 36370
rect 28590 36318 28642 36370
rect 31950 36318 32002 36370
rect 11902 36206 11954 36258
rect 12798 36206 12850 36258
rect 16270 36206 16322 36258
rect 19630 36206 19682 36258
rect 20190 36206 20242 36258
rect 20414 36206 20466 36258
rect 21310 36206 21362 36258
rect 21534 36206 21586 36258
rect 22206 36206 22258 36258
rect 22542 36206 22594 36258
rect 26574 36206 26626 36258
rect 35758 36206 35810 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 11342 35870 11394 35922
rect 12238 35870 12290 35922
rect 13134 35870 13186 35922
rect 13582 35870 13634 35922
rect 14030 35870 14082 35922
rect 21422 35870 21474 35922
rect 21982 35870 22034 35922
rect 22206 35870 22258 35922
rect 22766 35870 22818 35922
rect 25342 35870 25394 35922
rect 25678 35870 25730 35922
rect 26238 35870 26290 35922
rect 26574 35870 26626 35922
rect 28366 35870 28418 35922
rect 28926 35870 28978 35922
rect 29374 35870 29426 35922
rect 29822 35870 29874 35922
rect 30718 35870 30770 35922
rect 30830 35870 30882 35922
rect 31950 35870 32002 35922
rect 33182 35870 33234 35922
rect 34414 35870 34466 35922
rect 12014 35758 12066 35810
rect 13918 35758 13970 35810
rect 14478 35758 14530 35810
rect 14926 35758 14978 35810
rect 15150 35758 15202 35810
rect 15710 35758 15762 35810
rect 15934 35758 15986 35810
rect 16382 35758 16434 35810
rect 19630 35758 19682 35810
rect 23550 35758 23602 35810
rect 23662 35758 23714 35810
rect 24670 35758 24722 35810
rect 27134 35758 27186 35810
rect 11006 35646 11058 35698
rect 11230 35646 11282 35698
rect 11454 35646 11506 35698
rect 11902 35646 11954 35698
rect 12350 35646 12402 35698
rect 14366 35646 14418 35698
rect 14702 35646 14754 35698
rect 16270 35646 16322 35698
rect 16494 35646 16546 35698
rect 16942 35646 16994 35698
rect 17838 35646 17890 35698
rect 19182 35646 19234 35698
rect 19742 35646 19794 35698
rect 21086 35646 21138 35698
rect 21310 35646 21362 35698
rect 21534 35646 21586 35698
rect 21758 35646 21810 35698
rect 22318 35646 22370 35698
rect 22654 35646 22706 35698
rect 23886 35646 23938 35698
rect 24222 35646 24274 35698
rect 25230 35646 25282 35698
rect 25454 35646 25506 35698
rect 26686 35646 26738 35698
rect 27358 35646 27410 35698
rect 30606 35646 30658 35698
rect 31166 35646 31218 35698
rect 31838 35646 31890 35698
rect 32062 35646 32114 35698
rect 32510 35646 32562 35698
rect 32958 35646 33010 35698
rect 33294 35646 33346 35698
rect 33742 35646 33794 35698
rect 9998 35534 10050 35586
rect 10558 35534 10610 35586
rect 15150 35534 15202 35586
rect 15710 35534 15762 35586
rect 17390 35534 17442 35586
rect 18174 35534 18226 35586
rect 18734 35534 18786 35586
rect 20302 35534 20354 35586
rect 20750 35534 20802 35586
rect 27918 35534 27970 35586
rect 28814 35534 28866 35586
rect 30270 35534 30322 35586
rect 34302 35534 34354 35586
rect 34862 35534 34914 35586
rect 22766 35422 22818 35474
rect 23998 35422 24050 35474
rect 24334 35422 24386 35474
rect 24558 35422 24610 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 7310 35086 7362 35138
rect 7982 35086 8034 35138
rect 15486 35086 15538 35138
rect 20750 35086 20802 35138
rect 25454 35086 25506 35138
rect 26126 35086 26178 35138
rect 7534 34974 7586 35026
rect 7982 34974 8034 35026
rect 8654 34974 8706 35026
rect 10558 34974 10610 35026
rect 12462 34974 12514 35026
rect 14814 34974 14866 35026
rect 16270 34974 16322 35026
rect 19406 34974 19458 35026
rect 19854 34974 19906 35026
rect 20414 34974 20466 35026
rect 20638 34974 20690 35026
rect 22990 34974 23042 35026
rect 24558 34974 24610 35026
rect 29710 34974 29762 35026
rect 30270 34974 30322 35026
rect 31838 34974 31890 35026
rect 32510 34974 32562 35026
rect 33406 34974 33458 35026
rect 7086 34862 7138 34914
rect 8766 34862 8818 34914
rect 9774 34862 9826 34914
rect 10670 34862 10722 34914
rect 11678 34862 11730 34914
rect 11902 34862 11954 34914
rect 14030 34862 14082 34914
rect 14478 34862 14530 34914
rect 16046 34862 16098 34914
rect 16494 34862 16546 34914
rect 16830 34862 16882 34914
rect 17502 34862 17554 34914
rect 17726 34862 17778 34914
rect 18062 34862 18114 34914
rect 18398 34862 18450 34914
rect 22206 34862 22258 34914
rect 22430 34862 22482 34914
rect 23214 34862 23266 34914
rect 23438 34862 23490 34914
rect 24222 34862 24274 34914
rect 25678 34862 25730 34914
rect 27134 34862 27186 34914
rect 31390 34862 31442 34914
rect 32062 34862 32114 34914
rect 33966 34862 34018 34914
rect 9998 34750 10050 34802
rect 11006 34750 11058 34802
rect 13918 34750 13970 34802
rect 14142 34750 14194 34802
rect 15822 34750 15874 34802
rect 18286 34750 18338 34802
rect 18846 34750 18898 34802
rect 18958 34750 19010 34802
rect 22654 34750 22706 34802
rect 24558 34750 24610 34802
rect 25230 34750 25282 34802
rect 26574 34750 26626 34802
rect 26910 34750 26962 34802
rect 28142 34750 28194 34802
rect 28254 34750 28306 34802
rect 32398 34750 32450 34802
rect 32734 34750 32786 34802
rect 32958 34750 33010 34802
rect 6750 34638 6802 34690
rect 6974 34638 7026 34690
rect 9102 34638 9154 34690
rect 9214 34638 9266 34690
rect 9326 34638 9378 34690
rect 10222 34638 10274 34690
rect 10446 34638 10498 34690
rect 13022 34638 13074 34690
rect 14702 34638 14754 34690
rect 15262 34638 15314 34690
rect 15374 34638 15426 34690
rect 16270 34638 16322 34690
rect 18622 34638 18674 34690
rect 23886 34638 23938 34690
rect 24334 34638 24386 34690
rect 24670 34638 24722 34690
rect 26126 34638 26178 34690
rect 27246 34638 27298 34690
rect 27358 34638 27410 34690
rect 27470 34638 27522 34690
rect 27918 34638 27970 34690
rect 29374 34638 29426 34690
rect 30942 34638 30994 34690
rect 31614 34638 31666 34690
rect 31838 34638 31890 34690
rect 33518 34638 33570 34690
rect 34414 34638 34466 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 7422 34302 7474 34354
rect 14478 34302 14530 34354
rect 14702 34302 14754 34354
rect 14926 34302 14978 34354
rect 16942 34302 16994 34354
rect 17502 34302 17554 34354
rect 18510 34302 18562 34354
rect 18734 34302 18786 34354
rect 25454 34302 25506 34354
rect 29374 34302 29426 34354
rect 30718 34302 30770 34354
rect 30830 34302 30882 34354
rect 6638 34190 6690 34242
rect 11342 34190 11394 34242
rect 13918 34190 13970 34242
rect 16718 34190 16770 34242
rect 21086 34190 21138 34242
rect 21422 34190 21474 34242
rect 25678 34190 25730 34242
rect 27582 34190 27634 34242
rect 27918 34190 27970 34242
rect 31390 34190 31442 34242
rect 3950 34078 4002 34130
rect 4286 34078 4338 34130
rect 8542 34078 8594 34130
rect 8878 34078 8930 34130
rect 10110 34078 10162 34130
rect 10782 34078 10834 34130
rect 11454 34078 11506 34130
rect 12014 34078 12066 34130
rect 12686 34078 12738 34130
rect 14030 34078 14082 34130
rect 15374 34078 15426 34130
rect 15598 34078 15650 34130
rect 16606 34078 16658 34130
rect 17390 34078 17442 34130
rect 17614 34078 17666 34130
rect 19182 34078 19234 34130
rect 20638 34078 20690 34130
rect 20974 34078 21026 34130
rect 22094 34078 22146 34130
rect 22318 34078 22370 34130
rect 23326 34078 23378 34130
rect 24110 34078 24162 34130
rect 24334 34078 24386 34130
rect 24670 34078 24722 34130
rect 25230 34078 25282 34130
rect 26238 34078 26290 34130
rect 27134 34078 27186 34130
rect 27358 34078 27410 34130
rect 28030 34078 28082 34130
rect 28478 34078 28530 34130
rect 30494 34078 30546 34130
rect 30606 34078 30658 34130
rect 31054 34078 31106 34130
rect 32286 34078 32338 34130
rect 33630 34078 33682 34130
rect 8990 33966 9042 34018
rect 12798 33966 12850 34018
rect 14814 33966 14866 34018
rect 16270 33966 16322 34018
rect 18622 33966 18674 34018
rect 19518 33966 19570 34018
rect 23438 33966 23490 34018
rect 23774 33966 23826 34018
rect 24222 33966 24274 34018
rect 25342 33966 25394 34018
rect 26126 33966 26178 34018
rect 29822 33966 29874 34018
rect 32174 33966 32226 34018
rect 33294 33966 33346 34018
rect 34078 33966 34130 34018
rect 10222 33854 10274 33906
rect 13918 33854 13970 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 6974 33518 7026 33570
rect 10558 33518 10610 33570
rect 12126 33518 12178 33570
rect 14590 33518 14642 33570
rect 24558 33518 24610 33570
rect 27918 33518 27970 33570
rect 6190 33406 6242 33458
rect 8094 33406 8146 33458
rect 9998 33406 10050 33458
rect 15038 33406 15090 33458
rect 15822 33406 15874 33458
rect 16494 33406 16546 33458
rect 19070 33406 19122 33458
rect 23662 33406 23714 33458
rect 26126 33406 26178 33458
rect 27134 33406 27186 33458
rect 27582 33406 27634 33458
rect 28254 33406 28306 33458
rect 31614 33406 31666 33458
rect 31950 33406 32002 33458
rect 33630 33406 33682 33458
rect 6638 33294 6690 33346
rect 7870 33294 7922 33346
rect 8878 33294 8930 33346
rect 9662 33294 9714 33346
rect 10894 33294 10946 33346
rect 11454 33294 11506 33346
rect 11678 33294 11730 33346
rect 14702 33294 14754 33346
rect 15486 33294 15538 33346
rect 16382 33294 16434 33346
rect 16606 33294 16658 33346
rect 17054 33294 17106 33346
rect 17614 33294 17666 33346
rect 18846 33294 18898 33346
rect 21758 33294 21810 33346
rect 21982 33294 22034 33346
rect 22430 33294 22482 33346
rect 23214 33294 23266 33346
rect 23550 33294 23602 33346
rect 23998 33294 24050 33346
rect 24222 33294 24274 33346
rect 25118 33294 25170 33346
rect 26910 33294 26962 33346
rect 30382 33294 30434 33346
rect 31502 33294 31554 33346
rect 32734 33294 32786 33346
rect 33182 33294 33234 33346
rect 33742 33294 33794 33346
rect 34190 33294 34242 33346
rect 35086 33294 35138 33346
rect 35310 33294 35362 33346
rect 7086 33182 7138 33234
rect 8542 33182 8594 33234
rect 9102 33182 9154 33234
rect 11118 33182 11170 33234
rect 17838 33182 17890 33234
rect 18398 33182 18450 33234
rect 18734 33182 18786 33234
rect 21870 33182 21922 33234
rect 25006 33182 25058 33234
rect 28142 33182 28194 33234
rect 30494 33182 30546 33234
rect 32286 33182 32338 33234
rect 34974 33182 35026 33234
rect 6078 33070 6130 33122
rect 6302 33070 6354 33122
rect 8206 33070 8258 33122
rect 8654 33070 8706 33122
rect 9550 33070 9602 33122
rect 19182 33070 19234 33122
rect 19406 33070 19458 33122
rect 19966 33070 20018 33122
rect 24782 33070 24834 33122
rect 26238 33070 26290 33122
rect 30718 33070 30770 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 13582 32734 13634 32786
rect 15150 32734 15202 32786
rect 16830 32734 16882 32786
rect 23326 32734 23378 32786
rect 27134 32734 27186 32786
rect 30830 32734 30882 32786
rect 33406 32734 33458 32786
rect 8654 32622 8706 32674
rect 9998 32622 10050 32674
rect 10446 32622 10498 32674
rect 10894 32622 10946 32674
rect 12574 32622 12626 32674
rect 13694 32622 13746 32674
rect 18286 32622 18338 32674
rect 19294 32622 19346 32674
rect 22654 32622 22706 32674
rect 24110 32622 24162 32674
rect 26910 32622 26962 32674
rect 27918 32622 27970 32674
rect 28030 32622 28082 32674
rect 30606 32622 30658 32674
rect 31054 32622 31106 32674
rect 34078 32622 34130 32674
rect 8206 32510 8258 32562
rect 9886 32510 9938 32562
rect 10110 32510 10162 32562
rect 10670 32510 10722 32562
rect 11006 32510 11058 32562
rect 12798 32510 12850 32562
rect 14702 32510 14754 32562
rect 14926 32510 14978 32562
rect 17726 32510 17778 32562
rect 19406 32510 19458 32562
rect 22766 32510 22818 32562
rect 23214 32510 23266 32562
rect 23550 32510 23602 32562
rect 23998 32510 24050 32562
rect 24222 32510 24274 32562
rect 24670 32510 24722 32562
rect 27246 32510 27298 32562
rect 27358 32510 27410 32562
rect 30494 32510 30546 32562
rect 31726 32510 31778 32562
rect 32958 32510 33010 32562
rect 33630 32510 33682 32562
rect 33854 32510 33906 32562
rect 34190 32510 34242 32562
rect 6078 32398 6130 32450
rect 6862 32398 6914 32450
rect 7310 32398 7362 32450
rect 7758 32398 7810 32450
rect 11454 32398 11506 32450
rect 14142 32398 14194 32450
rect 14814 32398 14866 32450
rect 16382 32398 16434 32450
rect 20974 32398 21026 32450
rect 31390 32398 31442 32450
rect 33518 32398 33570 32450
rect 13134 32286 13186 32338
rect 13582 32286 13634 32338
rect 14030 32286 14082 32338
rect 27918 32286 27970 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 7758 31950 7810 32002
rect 5854 31838 5906 31890
rect 6302 31838 6354 31890
rect 6862 31838 6914 31890
rect 19406 31838 19458 31890
rect 24222 31838 24274 31890
rect 26350 31838 26402 31890
rect 28030 31838 28082 31890
rect 28478 31838 28530 31890
rect 30942 31838 30994 31890
rect 33182 31838 33234 31890
rect 7758 31726 7810 31778
rect 13582 31726 13634 31778
rect 15262 31726 15314 31778
rect 17278 31726 17330 31778
rect 18622 31726 18674 31778
rect 22206 31726 22258 31778
rect 22430 31726 22482 31778
rect 23438 31726 23490 31778
rect 23886 31726 23938 31778
rect 24446 31726 24498 31778
rect 25678 31726 25730 31778
rect 26574 31726 26626 31778
rect 27022 31726 27074 31778
rect 27918 31726 27970 31778
rect 28142 31726 28194 31778
rect 29150 31726 29202 31778
rect 31278 31726 31330 31778
rect 31838 31726 31890 31778
rect 32062 31726 32114 31778
rect 32510 31726 32562 31778
rect 33742 31726 33794 31778
rect 2046 31614 2098 31666
rect 7310 31614 7362 31666
rect 8094 31614 8146 31666
rect 8878 31614 8930 31666
rect 9214 31614 9266 31666
rect 11454 31614 11506 31666
rect 11566 31614 11618 31666
rect 13470 31614 13522 31666
rect 15598 31614 15650 31666
rect 17054 31614 17106 31666
rect 18398 31614 18450 31666
rect 19294 31614 19346 31666
rect 23214 31614 23266 31666
rect 24110 31614 24162 31666
rect 26014 31614 26066 31666
rect 26910 31614 26962 31666
rect 27582 31614 27634 31666
rect 28590 31614 28642 31666
rect 29262 31614 29314 31666
rect 29822 31614 29874 31666
rect 30606 31614 30658 31666
rect 30830 31614 30882 31666
rect 31502 31614 31554 31666
rect 32734 31614 32786 31666
rect 33406 31614 33458 31666
rect 33854 31614 33906 31666
rect 39566 31614 39618 31666
rect 1710 31502 1762 31554
rect 2494 31502 2546 31554
rect 5742 31502 5794 31554
rect 7422 31502 7474 31554
rect 8542 31502 8594 31554
rect 8766 31502 8818 31554
rect 9326 31502 9378 31554
rect 9550 31502 9602 31554
rect 11790 31502 11842 31554
rect 18734 31502 18786 31554
rect 18846 31502 18898 31554
rect 22766 31502 22818 31554
rect 23326 31502 23378 31554
rect 25902 31502 25954 31554
rect 26798 31502 26850 31554
rect 31726 31502 31778 31554
rect 32286 31502 32338 31554
rect 34078 31502 34130 31554
rect 39230 31502 39282 31554
rect 39902 31502 39954 31554
rect 40238 31502 40290 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 3278 31166 3330 31218
rect 10558 31166 10610 31218
rect 11118 31166 11170 31218
rect 14702 31166 14754 31218
rect 15374 31166 15426 31218
rect 15598 31166 15650 31218
rect 16718 31166 16770 31218
rect 19518 31166 19570 31218
rect 20750 31166 20802 31218
rect 26126 31166 26178 31218
rect 31614 31166 31666 31218
rect 33070 31166 33122 31218
rect 39902 31166 39954 31218
rect 6526 31054 6578 31106
rect 6638 31054 6690 31106
rect 8542 31054 8594 31106
rect 8766 31054 8818 31106
rect 9550 31054 9602 31106
rect 13470 31054 13522 31106
rect 13806 31054 13858 31106
rect 16606 31054 16658 31106
rect 16830 31054 16882 31106
rect 18510 31054 18562 31106
rect 20638 31054 20690 31106
rect 31502 31054 31554 31106
rect 33294 31054 33346 31106
rect 5630 30942 5682 30994
rect 6190 30942 6242 30994
rect 7758 30942 7810 30994
rect 8094 30942 8146 30994
rect 9662 30942 9714 30994
rect 9886 30942 9938 30994
rect 10110 30942 10162 30994
rect 11006 30942 11058 30994
rect 11342 30942 11394 30994
rect 11454 30942 11506 30994
rect 12126 30942 12178 30994
rect 13022 30942 13074 30994
rect 13918 30942 13970 30994
rect 15038 30942 15090 30994
rect 15486 30942 15538 30994
rect 17502 30942 17554 30994
rect 17950 30942 18002 30994
rect 18174 30942 18226 30994
rect 18734 30942 18786 30994
rect 18958 30942 19010 30994
rect 19406 30942 19458 30994
rect 19966 30942 20018 30994
rect 20974 30942 21026 30994
rect 22878 30942 22930 30994
rect 26014 30942 26066 30994
rect 26798 30942 26850 30994
rect 28478 30942 28530 30994
rect 32174 30942 32226 30994
rect 32398 30942 32450 30994
rect 33742 30942 33794 30994
rect 40238 30942 40290 30994
rect 7198 30830 7250 30882
rect 8878 30830 8930 30882
rect 14254 30830 14306 30882
rect 14590 30830 14642 30882
rect 17726 30830 17778 30882
rect 19182 30830 19234 30882
rect 19742 30830 19794 30882
rect 22542 30830 22594 30882
rect 23326 30830 23378 30882
rect 27022 30830 27074 30882
rect 27470 30830 27522 30882
rect 27806 30830 27858 30882
rect 28254 30830 28306 30882
rect 30718 30830 30770 30882
rect 31278 30830 31330 30882
rect 32062 30830 32114 30882
rect 33182 30830 33234 30882
rect 2494 30718 2546 30770
rect 6526 30718 6578 30770
rect 20302 30718 20354 30770
rect 32510 30718 32562 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 14254 30382 14306 30434
rect 18286 30382 18338 30434
rect 21310 30382 21362 30434
rect 26126 30382 26178 30434
rect 8094 30270 8146 30322
rect 9774 30270 9826 30322
rect 10446 30270 10498 30322
rect 14030 30270 14082 30322
rect 15374 30270 15426 30322
rect 17390 30270 17442 30322
rect 18174 30270 18226 30322
rect 19406 30270 19458 30322
rect 21422 30270 21474 30322
rect 2158 30158 2210 30210
rect 2830 30158 2882 30210
rect 6078 30158 6130 30210
rect 6750 30158 6802 30210
rect 6974 30158 7026 30210
rect 8206 30158 8258 30210
rect 8878 30158 8930 30210
rect 9326 30158 9378 30210
rect 10222 30158 10274 30210
rect 11902 30158 11954 30210
rect 12238 30158 12290 30210
rect 12462 30158 12514 30210
rect 12798 30158 12850 30210
rect 13806 30158 13858 30210
rect 14478 30158 14530 30210
rect 15486 30158 15538 30210
rect 17166 30158 17218 30210
rect 17950 30158 18002 30210
rect 18622 30158 18674 30210
rect 19182 30158 19234 30210
rect 20078 30158 20130 30210
rect 20526 30158 20578 30210
rect 21646 30158 21698 30210
rect 22766 30158 22818 30210
rect 23326 30158 23378 30210
rect 27470 30158 27522 30210
rect 27918 30158 27970 30210
rect 29150 30158 29202 30210
rect 29262 30158 29314 30210
rect 30942 30158 30994 30210
rect 31278 30158 31330 30210
rect 33518 30158 33570 30210
rect 35646 30158 35698 30210
rect 6302 30046 6354 30098
rect 6526 30046 6578 30098
rect 7310 30046 7362 30098
rect 9438 30046 9490 30098
rect 10558 30046 10610 30098
rect 12014 30046 12066 30098
rect 12574 30046 12626 30098
rect 16158 30046 16210 30098
rect 17614 30046 17666 30098
rect 20414 30046 20466 30098
rect 24222 30046 24274 30098
rect 25006 30046 25058 30098
rect 26350 30046 26402 30098
rect 26910 30046 26962 30098
rect 27358 30046 27410 30098
rect 30606 30046 30658 30098
rect 31950 30046 32002 30098
rect 34974 30046 35026 30098
rect 5182 29934 5234 29986
rect 6638 29934 6690 29986
rect 14926 29934 14978 29986
rect 20190 29934 20242 29986
rect 20302 29934 20354 29986
rect 22094 29934 22146 29986
rect 25454 29934 25506 29986
rect 25790 29934 25842 29986
rect 29822 29934 29874 29986
rect 30382 29934 30434 29986
rect 31054 29934 31106 29986
rect 33966 29934 34018 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 5742 29598 5794 29650
rect 7086 29598 7138 29650
rect 9102 29598 9154 29650
rect 10222 29598 10274 29650
rect 10446 29598 10498 29650
rect 10894 29598 10946 29650
rect 14590 29598 14642 29650
rect 17614 29598 17666 29650
rect 19406 29598 19458 29650
rect 20414 29598 20466 29650
rect 32062 29598 32114 29650
rect 32510 29598 32562 29650
rect 34526 29598 34578 29650
rect 2046 29486 2098 29538
rect 8430 29486 8482 29538
rect 8766 29486 8818 29538
rect 8878 29486 8930 29538
rect 9886 29486 9938 29538
rect 13694 29486 13746 29538
rect 15486 29486 15538 29538
rect 17502 29486 17554 29538
rect 19070 29486 19122 29538
rect 24334 29486 24386 29538
rect 24670 29486 24722 29538
rect 31390 29486 31442 29538
rect 1710 29374 1762 29426
rect 5630 29374 5682 29426
rect 5854 29374 5906 29426
rect 6190 29374 6242 29426
rect 7534 29374 7586 29426
rect 7982 29374 8034 29426
rect 9774 29374 9826 29426
rect 10110 29374 10162 29426
rect 10558 29374 10610 29426
rect 13582 29374 13634 29426
rect 14702 29374 14754 29426
rect 16158 29374 16210 29426
rect 16382 29374 16434 29426
rect 18174 29374 18226 29426
rect 18622 29374 18674 29426
rect 19518 29374 19570 29426
rect 19630 29374 19682 29426
rect 20078 29374 20130 29426
rect 20302 29374 20354 29426
rect 26350 29374 26402 29426
rect 33518 29374 33570 29426
rect 33966 29374 34018 29426
rect 34750 29374 34802 29426
rect 35198 29374 35250 29426
rect 35422 29374 35474 29426
rect 39006 29374 39058 29426
rect 2494 29262 2546 29314
rect 5294 29262 5346 29314
rect 6190 29262 6242 29314
rect 6414 29262 6466 29314
rect 6638 29262 6690 29314
rect 11006 29262 11058 29314
rect 20974 29262 21026 29314
rect 25230 29262 25282 29314
rect 25790 29262 25842 29314
rect 33070 29262 33122 29314
rect 34638 29262 34690 29314
rect 34974 29262 35026 29314
rect 35870 29262 35922 29314
rect 40126 29262 40178 29314
rect 17614 29150 17666 29202
rect 20414 29150 20466 29202
rect 25342 29150 25394 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 11790 28814 11842 28866
rect 12910 28814 12962 28866
rect 16718 28814 16770 28866
rect 17838 28814 17890 28866
rect 26686 28814 26738 28866
rect 31054 28814 31106 28866
rect 32510 28814 32562 28866
rect 8318 28702 8370 28754
rect 9214 28702 9266 28754
rect 10110 28702 10162 28754
rect 11902 28702 11954 28754
rect 12910 28702 12962 28754
rect 14142 28702 14194 28754
rect 15486 28702 15538 28754
rect 16942 28702 16994 28754
rect 17950 28702 18002 28754
rect 19966 28702 20018 28754
rect 21422 28702 21474 28754
rect 21758 28702 21810 28754
rect 27358 28702 27410 28754
rect 27582 28702 27634 28754
rect 27918 28702 27970 28754
rect 28590 28702 28642 28754
rect 29598 28702 29650 28754
rect 31502 28702 31554 28754
rect 33966 28702 34018 28754
rect 35534 28702 35586 28754
rect 2942 28590 2994 28642
rect 6414 28590 6466 28642
rect 6638 28590 6690 28642
rect 6974 28590 7026 28642
rect 7646 28590 7698 28642
rect 8206 28590 8258 28642
rect 8990 28590 9042 28642
rect 10446 28590 10498 28642
rect 11454 28590 11506 28642
rect 12462 28590 12514 28642
rect 13582 28590 13634 28642
rect 15150 28590 15202 28642
rect 15934 28590 15986 28642
rect 17390 28590 17442 28642
rect 22654 28590 22706 28642
rect 22990 28590 23042 28642
rect 23662 28590 23714 28642
rect 29150 28590 29202 28642
rect 30382 28590 30434 28642
rect 31278 28590 31330 28642
rect 31726 28590 31778 28642
rect 31950 28590 32002 28642
rect 33518 28590 33570 28642
rect 34302 28590 34354 28642
rect 34750 28590 34802 28642
rect 35422 28590 35474 28642
rect 36318 28590 36370 28642
rect 37102 28590 37154 28642
rect 37550 28590 37602 28642
rect 39678 28590 39730 28642
rect 40238 28590 40290 28642
rect 6862 28478 6914 28530
rect 9662 28478 9714 28530
rect 11006 28478 11058 28530
rect 13694 28478 13746 28530
rect 16270 28478 16322 28530
rect 17278 28478 17330 28530
rect 25902 28478 25954 28530
rect 27022 28478 27074 28530
rect 27806 28478 27858 28530
rect 28030 28478 28082 28530
rect 32398 28478 32450 28530
rect 32510 28478 32562 28530
rect 33406 28478 33458 28530
rect 39902 28478 39954 28530
rect 2158 28366 2210 28418
rect 5854 28366 5906 28418
rect 5966 28366 6018 28418
rect 6078 28366 6130 28418
rect 17166 28366 17218 28418
rect 18398 28366 18450 28418
rect 19070 28366 19122 28418
rect 21870 28366 21922 28418
rect 31838 28366 31890 28418
rect 36094 28366 36146 28418
rect 36990 28366 37042 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 6750 28030 6802 28082
rect 7310 28030 7362 28082
rect 7534 28030 7586 28082
rect 8766 28030 8818 28082
rect 10334 28030 10386 28082
rect 10446 28030 10498 28082
rect 10558 28030 10610 28082
rect 14702 28030 14754 28082
rect 16606 28030 16658 28082
rect 17726 28030 17778 28082
rect 21758 28030 21810 28082
rect 22542 28030 22594 28082
rect 22766 28030 22818 28082
rect 23774 28030 23826 28082
rect 24334 28030 24386 28082
rect 26350 28030 26402 28082
rect 29710 28030 29762 28082
rect 30718 28030 30770 28082
rect 32958 28030 33010 28082
rect 33182 28030 33234 28082
rect 36878 28030 36930 28082
rect 37438 28030 37490 28082
rect 8654 27918 8706 27970
rect 23550 27918 23602 27970
rect 23886 27918 23938 27970
rect 30830 27918 30882 27970
rect 33294 27918 33346 27970
rect 3838 27806 3890 27858
rect 4286 27806 4338 27858
rect 10222 27806 10274 27858
rect 10782 27806 10834 27858
rect 11790 27806 11842 27858
rect 12238 27806 12290 27858
rect 19070 27806 19122 27858
rect 19518 27806 19570 27858
rect 22990 27806 23042 27858
rect 23438 27806 23490 27858
rect 26574 27806 26626 27858
rect 27246 27806 27298 27858
rect 30382 27806 30434 27858
rect 31950 27806 32002 27858
rect 33742 27806 33794 27858
rect 34414 27806 34466 27858
rect 7646 27694 7698 27746
rect 8094 27694 8146 27746
rect 11454 27694 11506 27746
rect 15934 27694 15986 27746
rect 22878 27694 22930 27746
rect 25342 27694 25394 27746
rect 31502 27694 31554 27746
rect 32286 27694 32338 27746
rect 15374 27582 15426 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 10446 27246 10498 27298
rect 17054 27246 17106 27298
rect 29598 27246 29650 27298
rect 30718 27246 30770 27298
rect 31502 27246 31554 27298
rect 31726 27246 31778 27298
rect 33854 27246 33906 27298
rect 35198 27246 35250 27298
rect 7422 27134 7474 27186
rect 10782 27134 10834 27186
rect 12238 27134 12290 27186
rect 25454 27134 25506 27186
rect 26686 27134 26738 27186
rect 27470 27134 27522 27186
rect 28590 27134 28642 27186
rect 33406 27134 33458 27186
rect 33854 27134 33906 27186
rect 34750 27134 34802 27186
rect 35198 27134 35250 27186
rect 13358 27022 13410 27074
rect 14030 27022 14082 27074
rect 18286 27022 18338 27074
rect 19406 27022 19458 27074
rect 21198 27022 21250 27074
rect 21870 27022 21922 27074
rect 25006 27022 25058 27074
rect 25902 27022 25954 27074
rect 26238 27022 26290 27074
rect 30942 27022 30994 27074
rect 32174 27022 32226 27074
rect 32510 27022 32562 27074
rect 8430 26910 8482 26962
rect 10670 26910 10722 26962
rect 11118 26910 11170 26962
rect 11230 26910 11282 26962
rect 12350 26910 12402 26962
rect 17390 26910 17442 26962
rect 27806 26910 27858 26962
rect 28142 26910 28194 26962
rect 29262 26910 29314 26962
rect 29822 26910 29874 26962
rect 30382 26910 30434 26962
rect 32286 26910 32338 26962
rect 10222 26798 10274 26850
rect 11342 26798 11394 26850
rect 12126 26798 12178 26850
rect 12574 26798 12626 26850
rect 16270 26798 16322 26850
rect 18958 26798 19010 26850
rect 24110 26798 24162 26850
rect 31390 26798 31442 26850
rect 33070 26798 33122 26850
rect 34302 26798 34354 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 6414 26462 6466 26514
rect 7758 26462 7810 26514
rect 16046 26462 16098 26514
rect 23102 26462 23154 26514
rect 23886 26462 23938 26514
rect 33406 26462 33458 26514
rect 34414 26462 34466 26514
rect 7534 26350 7586 26402
rect 8654 26350 8706 26402
rect 13358 26350 13410 26402
rect 23214 26350 23266 26402
rect 31950 26350 32002 26402
rect 32510 26350 32562 26402
rect 2830 26238 2882 26290
rect 7982 26238 8034 26290
rect 8094 26238 8146 26290
rect 8542 26238 8594 26290
rect 8878 26238 8930 26290
rect 9662 26238 9714 26290
rect 15486 26238 15538 26290
rect 15934 26238 15986 26290
rect 16494 26238 16546 26290
rect 18510 26238 18562 26290
rect 19966 26238 20018 26290
rect 21982 26238 22034 26290
rect 22430 26238 22482 26290
rect 22766 26238 22818 26290
rect 22990 26238 23042 26290
rect 23438 26238 23490 26290
rect 26350 26238 26402 26290
rect 26686 26238 26738 26290
rect 29038 26238 29090 26290
rect 29486 26238 29538 26290
rect 29710 26238 29762 26290
rect 31166 26238 31218 26290
rect 32174 26238 32226 26290
rect 32958 26238 33010 26290
rect 33294 26238 33346 26290
rect 33966 26238 34018 26290
rect 39006 26238 39058 26290
rect 1934 26126 1986 26178
rect 6974 26126 7026 26178
rect 7870 26126 7922 26178
rect 17950 26126 18002 26178
rect 18622 26126 18674 26178
rect 19070 26126 19122 26178
rect 19294 26126 19346 26178
rect 21534 26126 21586 26178
rect 23774 26126 23826 26178
rect 24334 26126 24386 26178
rect 27358 26126 27410 26178
rect 28478 26126 28530 26178
rect 28814 26126 28866 26178
rect 29262 26126 29314 26178
rect 30382 26126 30434 26178
rect 30718 26126 30770 26178
rect 31614 26126 31666 26178
rect 32062 26126 32114 26178
rect 33742 26126 33794 26178
rect 34862 26126 34914 26178
rect 35310 26126 35362 26178
rect 40126 26126 40178 26178
rect 19406 26014 19458 26066
rect 33518 26014 33570 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 8766 25678 8818 25730
rect 13582 25678 13634 25730
rect 14702 25678 14754 25730
rect 20302 25678 20354 25730
rect 21534 25678 21586 25730
rect 36542 25678 36594 25730
rect 7310 25566 7362 25618
rect 10446 25566 10498 25618
rect 12126 25566 12178 25618
rect 12574 25566 12626 25618
rect 12686 25566 12738 25618
rect 14814 25566 14866 25618
rect 15262 25566 15314 25618
rect 16382 25566 16434 25618
rect 23774 25566 23826 25618
rect 24222 25566 24274 25618
rect 2942 25454 2994 25506
rect 4734 25454 4786 25506
rect 5070 25454 5122 25506
rect 5630 25454 5682 25506
rect 5854 25454 5906 25506
rect 6190 25454 6242 25506
rect 6414 25454 6466 25506
rect 6750 25454 6802 25506
rect 7982 25454 8034 25506
rect 8206 25454 8258 25506
rect 9438 25454 9490 25506
rect 9774 25454 9826 25506
rect 10334 25454 10386 25506
rect 11566 25454 11618 25506
rect 12014 25454 12066 25506
rect 13694 25454 13746 25506
rect 14366 25454 14418 25506
rect 16606 25454 16658 25506
rect 17278 25454 17330 25506
rect 22430 25454 22482 25506
rect 22878 25454 22930 25506
rect 24782 25454 24834 25506
rect 25230 25454 25282 25506
rect 29598 25454 29650 25506
rect 29822 25454 29874 25506
rect 30046 25454 30098 25506
rect 30830 25454 30882 25506
rect 31502 25454 31554 25506
rect 32846 25454 32898 25506
rect 33406 25454 33458 25506
rect 39006 25454 39058 25506
rect 8654 25342 8706 25394
rect 9550 25342 9602 25394
rect 11230 25342 11282 25394
rect 12126 25342 12178 25394
rect 13582 25342 13634 25394
rect 14030 25342 14082 25394
rect 19518 25342 19570 25394
rect 21422 25342 21474 25394
rect 23326 25342 23378 25394
rect 30270 25342 30322 25394
rect 31726 25342 31778 25394
rect 2158 25230 2210 25282
rect 4958 25230 5010 25282
rect 5742 25230 5794 25282
rect 6638 25230 6690 25282
rect 8766 25230 8818 25282
rect 11790 25230 11842 25282
rect 12798 25230 12850 25282
rect 15710 25230 15762 25282
rect 20638 25230 20690 25282
rect 21534 25230 21586 25282
rect 27470 25230 27522 25282
rect 28254 25230 28306 25282
rect 28590 25230 28642 25282
rect 29822 25230 29874 25282
rect 32062 25230 32114 25282
rect 32174 25230 32226 25282
rect 32286 25230 32338 25282
rect 32510 25230 32562 25282
rect 35982 25230 36034 25282
rect 39790 25230 39842 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 2046 24894 2098 24946
rect 2830 24894 2882 24946
rect 3614 24894 3666 24946
rect 6862 24894 6914 24946
rect 10110 24894 10162 24946
rect 10222 24894 10274 24946
rect 13806 24894 13858 24946
rect 15822 24894 15874 24946
rect 18734 24894 18786 24946
rect 18846 24894 18898 24946
rect 19630 24894 19682 24946
rect 20302 24894 20354 24946
rect 21198 24894 21250 24946
rect 24446 24894 24498 24946
rect 25454 24894 25506 24946
rect 25902 24894 25954 24946
rect 26686 24894 26738 24946
rect 26798 24894 26850 24946
rect 27358 24894 27410 24946
rect 35982 24894 36034 24946
rect 36654 24894 36706 24946
rect 7982 24782 8034 24834
rect 9550 24782 9602 24834
rect 10446 24782 10498 24834
rect 11342 24782 11394 24834
rect 15262 24782 15314 24834
rect 17502 24782 17554 24834
rect 19406 24782 19458 24834
rect 19742 24782 19794 24834
rect 20526 24782 20578 24834
rect 22654 24782 22706 24834
rect 22990 24782 23042 24834
rect 23774 24782 23826 24834
rect 25790 24782 25842 24834
rect 26126 24782 26178 24834
rect 27246 24782 27298 24834
rect 30494 24782 30546 24834
rect 31502 24782 31554 24834
rect 33070 24782 33122 24834
rect 33182 24782 33234 24834
rect 36206 24782 36258 24834
rect 1710 24670 1762 24722
rect 5854 24670 5906 24722
rect 6526 24670 6578 24722
rect 8430 24670 8482 24722
rect 9998 24670 10050 24722
rect 11230 24670 11282 24722
rect 12910 24670 12962 24722
rect 14926 24670 14978 24722
rect 17390 24670 17442 24722
rect 17726 24670 17778 24722
rect 18622 24670 18674 24722
rect 19294 24670 19346 24722
rect 20190 24670 20242 24722
rect 20750 24670 20802 24722
rect 21086 24670 21138 24722
rect 21310 24670 21362 24722
rect 22094 24670 22146 24722
rect 23326 24670 23378 24722
rect 23998 24670 24050 24722
rect 24334 24670 24386 24722
rect 26238 24670 26290 24722
rect 26910 24670 26962 24722
rect 27582 24670 27634 24722
rect 28254 24670 28306 24722
rect 31726 24670 31778 24722
rect 32174 24670 32226 24722
rect 34302 24670 34354 24722
rect 35646 24670 35698 24722
rect 36318 24670 36370 24722
rect 2494 24558 2546 24610
rect 8878 24558 8930 24610
rect 16382 24558 16434 24610
rect 16830 24558 16882 24610
rect 18062 24558 18114 24610
rect 22206 24558 22258 24610
rect 23214 24558 23266 24610
rect 23662 24558 23714 24610
rect 31278 24558 31330 24610
rect 34414 24558 34466 24610
rect 35422 24558 35474 24610
rect 36766 24558 36818 24610
rect 37214 24558 37266 24610
rect 9662 24446 9714 24498
rect 17950 24446 18002 24498
rect 24446 24446 24498 24498
rect 33182 24446 33234 24498
rect 34190 24446 34242 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 9214 24110 9266 24162
rect 28478 24110 28530 24162
rect 29598 24110 29650 24162
rect 7646 23998 7698 24050
rect 8542 23998 8594 24050
rect 9550 23998 9602 24050
rect 10670 23998 10722 24050
rect 13694 23998 13746 24050
rect 14478 23998 14530 24050
rect 19406 23998 19458 24050
rect 20302 23998 20354 24050
rect 21758 23998 21810 24050
rect 27134 23998 27186 24050
rect 29486 23998 29538 24050
rect 33966 23998 34018 24050
rect 40014 23998 40066 24050
rect 2270 23886 2322 23938
rect 7086 23886 7138 23938
rect 7198 23886 7250 23938
rect 8094 23886 8146 23938
rect 10334 23886 10386 23938
rect 10558 23886 10610 23938
rect 12014 23886 12066 23938
rect 12574 23886 12626 23938
rect 14702 23886 14754 23938
rect 15374 23886 15426 23938
rect 20078 23886 20130 23938
rect 22430 23886 22482 23938
rect 23998 23886 24050 23938
rect 25006 23886 25058 23938
rect 25902 23886 25954 23938
rect 28254 23886 28306 23938
rect 28366 23886 28418 23938
rect 30382 23886 30434 23938
rect 33070 23886 33122 23938
rect 33518 23886 33570 23938
rect 34190 23886 34242 23938
rect 34638 23886 34690 23938
rect 35422 23886 35474 23938
rect 35870 23886 35922 23938
rect 39006 23886 39058 23938
rect 9438 23774 9490 23826
rect 11118 23774 11170 23826
rect 13470 23774 13522 23826
rect 18734 23774 18786 23826
rect 20750 23774 20802 23826
rect 21310 23774 21362 23826
rect 22990 23774 23042 23826
rect 26798 23774 26850 23826
rect 30494 23774 30546 23826
rect 1710 23662 1762 23714
rect 2718 23662 2770 23714
rect 17838 23662 17890 23714
rect 18398 23662 18450 23714
rect 21534 23662 21586 23714
rect 21758 23662 21810 23714
rect 21870 23662 21922 23714
rect 23326 23662 23378 23714
rect 27022 23662 27074 23714
rect 27246 23662 27298 23714
rect 27358 23662 27410 23714
rect 31166 23662 31218 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 3390 23326 3442 23378
rect 5406 23326 5458 23378
rect 16270 23326 16322 23378
rect 18398 23326 18450 23378
rect 19630 23326 19682 23378
rect 20078 23326 20130 23378
rect 20974 23326 21026 23378
rect 21198 23326 21250 23378
rect 22990 23326 23042 23378
rect 27358 23326 27410 23378
rect 33294 23326 33346 23378
rect 34862 23326 34914 23378
rect 39006 23326 39058 23378
rect 7310 23214 7362 23266
rect 8654 23214 8706 23266
rect 9662 23214 9714 23266
rect 12126 23214 12178 23266
rect 17502 23214 17554 23266
rect 25230 23214 25282 23266
rect 26686 23214 26738 23266
rect 34078 23214 34130 23266
rect 34638 23214 34690 23266
rect 39230 23214 39282 23266
rect 39902 23214 39954 23266
rect 2830 23102 2882 23154
rect 8318 23102 8370 23154
rect 8766 23102 8818 23154
rect 9550 23102 9602 23154
rect 11566 23102 11618 23154
rect 16158 23102 16210 23154
rect 17390 23102 17442 23154
rect 17614 23102 17666 23154
rect 17950 23102 18002 23154
rect 20414 23102 20466 23154
rect 22094 23158 22146 23210
rect 20638 23102 20690 23154
rect 22430 23102 22482 23154
rect 22654 23102 22706 23154
rect 24222 23102 24274 23154
rect 24558 23102 24610 23154
rect 25454 23102 25506 23154
rect 25902 23102 25954 23154
rect 26462 23102 26514 23154
rect 26798 23102 26850 23154
rect 27918 23102 27970 23154
rect 28590 23102 28642 23154
rect 31390 23102 31442 23154
rect 32174 23102 32226 23154
rect 33182 23102 33234 23154
rect 33966 23102 34018 23154
rect 34526 23102 34578 23154
rect 39566 23102 39618 23154
rect 40238 23102 40290 23154
rect 1934 22990 1986 23042
rect 8430 22990 8482 23042
rect 11454 22990 11506 23042
rect 16830 22990 16882 23042
rect 19294 22990 19346 23042
rect 19966 22990 20018 23042
rect 21870 22990 21922 23042
rect 24670 22990 24722 23042
rect 26238 22990 26290 23042
rect 27694 22990 27746 23042
rect 28702 22990 28754 23042
rect 31166 22990 31218 23042
rect 38558 22990 38610 23042
rect 16270 22878 16322 22930
rect 21646 22878 21698 22930
rect 25902 22878 25954 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 9998 22542 10050 22594
rect 28590 22542 28642 22594
rect 29486 22542 29538 22594
rect 29710 22542 29762 22594
rect 29934 22542 29986 22594
rect 34414 22542 34466 22594
rect 4846 22430 4898 22482
rect 5742 22430 5794 22482
rect 6750 22430 6802 22482
rect 7198 22430 7250 22482
rect 7534 22430 7586 22482
rect 7982 22430 8034 22482
rect 8654 22430 8706 22482
rect 11454 22430 11506 22482
rect 16158 22430 16210 22482
rect 17390 22430 17442 22482
rect 21646 22430 21698 22482
rect 22206 22430 22258 22482
rect 23102 22430 23154 22482
rect 25678 22430 25730 22482
rect 27134 22430 27186 22482
rect 27918 22430 27970 22482
rect 30158 22430 30210 22482
rect 30606 22430 30658 22482
rect 31614 22430 31666 22482
rect 35870 22430 35922 22482
rect 40014 22430 40066 22482
rect 2830 22318 2882 22370
rect 3838 22318 3890 22370
rect 8318 22318 8370 22370
rect 9214 22318 9266 22370
rect 11230 22318 11282 22370
rect 12014 22318 12066 22370
rect 12686 22318 12738 22370
rect 15934 22318 15986 22370
rect 17054 22318 17106 22370
rect 17614 22318 17666 22370
rect 18062 22318 18114 22370
rect 23326 22318 23378 22370
rect 25790 22318 25842 22370
rect 26238 22318 26290 22370
rect 29038 22318 29090 22370
rect 32958 22318 33010 22370
rect 33182 22318 33234 22370
rect 34974 22318 35026 22370
rect 39118 22318 39170 22370
rect 1934 22206 1986 22258
rect 3278 22206 3330 22258
rect 6190 22206 6242 22258
rect 8094 22206 8146 22258
rect 9550 22206 9602 22258
rect 9886 22206 9938 22258
rect 12910 22206 12962 22258
rect 16606 22206 16658 22258
rect 17166 22206 17218 22258
rect 18622 22206 18674 22258
rect 21758 22206 21810 22258
rect 22430 22206 22482 22258
rect 28478 22206 28530 22258
rect 32286 22206 32338 22258
rect 33406 22206 33458 22258
rect 33854 22206 33906 22258
rect 33966 22206 34018 22258
rect 34526 22206 34578 22258
rect 35422 22206 35474 22258
rect 2158 22094 2210 22146
rect 4734 22094 4786 22146
rect 6302 22094 6354 22146
rect 7310 22094 7362 22146
rect 8766 22094 8818 22146
rect 8878 22094 8930 22146
rect 9438 22094 9490 22146
rect 10446 22094 10498 22146
rect 10894 22094 10946 22146
rect 11902 22094 11954 22146
rect 14142 22094 14194 22146
rect 14590 22094 14642 22146
rect 17390 22094 17442 22146
rect 18174 22094 18226 22146
rect 18398 22094 18450 22146
rect 18734 22094 18786 22146
rect 18958 22094 19010 22146
rect 19294 22094 19346 22146
rect 19742 22094 19794 22146
rect 20302 22094 20354 22146
rect 20750 22094 20802 22146
rect 21534 22094 21586 22146
rect 22206 22094 22258 22146
rect 27470 22094 27522 22146
rect 31054 22094 31106 22146
rect 33294 22094 33346 22146
rect 33630 22094 33682 22146
rect 34414 22094 34466 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 1598 21758 1650 21810
rect 2382 21758 2434 21810
rect 5630 21758 5682 21810
rect 8542 21758 8594 21810
rect 9550 21758 9602 21810
rect 12910 21758 12962 21810
rect 13694 21758 13746 21810
rect 14702 21758 14754 21810
rect 17502 21758 17554 21810
rect 17614 21758 17666 21810
rect 25342 21758 25394 21810
rect 30942 21758 30994 21810
rect 33742 21758 33794 21810
rect 37438 21758 37490 21810
rect 38222 21758 38274 21810
rect 5742 21646 5794 21698
rect 7758 21646 7810 21698
rect 8766 21646 8818 21698
rect 10110 21646 10162 21698
rect 10446 21646 10498 21698
rect 12574 21646 12626 21698
rect 14478 21646 14530 21698
rect 15822 21646 15874 21698
rect 24222 21646 24274 21698
rect 27582 21646 27634 21698
rect 27918 21646 27970 21698
rect 29262 21646 29314 21698
rect 32174 21646 32226 21698
rect 33854 21646 33906 21698
rect 38334 21646 38386 21698
rect 4734 21534 4786 21586
rect 5294 21534 5346 21586
rect 5406 21534 5458 21586
rect 6190 21534 6242 21586
rect 6526 21534 6578 21586
rect 8094 21534 8146 21586
rect 8318 21534 8370 21586
rect 9774 21534 9826 21586
rect 12350 21534 12402 21586
rect 13470 21534 13522 21586
rect 14366 21534 14418 21586
rect 15262 21534 15314 21586
rect 15934 21534 15986 21586
rect 16494 21534 16546 21586
rect 18510 21534 18562 21586
rect 24334 21534 24386 21586
rect 25678 21534 25730 21586
rect 26910 21534 26962 21586
rect 28366 21534 28418 21586
rect 29710 21534 29762 21586
rect 30158 21534 30210 21586
rect 30606 21534 30658 21586
rect 30830 21534 30882 21586
rect 31166 21534 31218 21586
rect 32510 21534 32562 21586
rect 33630 21534 33682 21586
rect 33966 21534 34018 21586
rect 34526 21534 34578 21586
rect 34862 21534 34914 21586
rect 39006 21534 39058 21586
rect 8206 21422 8258 21474
rect 10558 21422 10610 21474
rect 11006 21422 11058 21474
rect 15486 21422 15538 21474
rect 18286 21422 18338 21474
rect 22318 21422 22370 21474
rect 28814 21422 28866 21474
rect 31726 21422 31778 21474
rect 40126 21422 40178 21474
rect 14926 21310 14978 21362
rect 17726 21310 17778 21362
rect 24222 21310 24274 21362
rect 31838 21310 31890 21362
rect 32510 21310 32562 21362
rect 33070 21310 33122 21362
rect 33294 21310 33346 21362
rect 37998 21310 38050 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 11790 20974 11842 21026
rect 12686 20974 12738 21026
rect 14478 20974 14530 21026
rect 19070 20974 19122 21026
rect 19630 20974 19682 21026
rect 20638 20974 20690 21026
rect 27582 20974 27634 21026
rect 29262 20974 29314 21026
rect 31502 20974 31554 21026
rect 33070 20974 33122 21026
rect 33966 20974 34018 21026
rect 35422 20974 35474 21026
rect 3726 20862 3778 20914
rect 4622 20862 4674 20914
rect 6302 20862 6354 20914
rect 7982 20862 8034 20914
rect 18622 20862 18674 20914
rect 19294 20862 19346 20914
rect 20190 20862 20242 20914
rect 22878 20862 22930 20914
rect 24222 20862 24274 20914
rect 24670 20862 24722 20914
rect 25454 20862 25506 20914
rect 26686 20862 26738 20914
rect 29822 20862 29874 20914
rect 30942 20862 30994 20914
rect 31950 20862 32002 20914
rect 33630 20862 33682 20914
rect 35534 20862 35586 20914
rect 1710 20750 1762 20802
rect 4286 20750 4338 20802
rect 4510 20750 4562 20802
rect 5182 20750 5234 20802
rect 6190 20750 6242 20802
rect 6750 20750 6802 20802
rect 6974 20750 7026 20802
rect 8430 20750 8482 20802
rect 8878 20750 8930 20802
rect 9662 20750 9714 20802
rect 12126 20750 12178 20802
rect 12350 20750 12402 20802
rect 13470 20750 13522 20802
rect 13694 20750 13746 20802
rect 13918 20750 13970 20802
rect 15374 20750 15426 20802
rect 15710 20750 15762 20802
rect 16494 20750 16546 20802
rect 17054 20750 17106 20802
rect 17614 20750 17666 20802
rect 18062 20750 18114 20802
rect 20750 20750 20802 20802
rect 22654 20750 22706 20802
rect 23102 20750 23154 20802
rect 23326 20750 23378 20802
rect 23998 20750 24050 20802
rect 25790 20750 25842 20802
rect 27694 20750 27746 20802
rect 31166 20750 31218 20802
rect 32846 20750 32898 20802
rect 33742 20750 33794 20802
rect 34414 20750 34466 20802
rect 35086 20750 35138 20802
rect 35198 20750 35250 20802
rect 37886 20750 37938 20802
rect 2270 20638 2322 20690
rect 3166 20638 3218 20690
rect 4734 20638 4786 20690
rect 7422 20638 7474 20690
rect 9550 20638 9602 20690
rect 10222 20638 10274 20690
rect 10446 20638 10498 20690
rect 11678 20638 11730 20690
rect 14366 20638 14418 20690
rect 15822 20638 15874 20690
rect 17166 20638 17218 20690
rect 18846 20638 18898 20690
rect 19854 20638 19906 20690
rect 20638 20638 20690 20690
rect 21758 20638 21810 20690
rect 22094 20638 22146 20690
rect 27358 20638 27410 20690
rect 29150 20638 29202 20690
rect 40238 20638 40290 20690
rect 2606 20526 2658 20578
rect 5966 20526 6018 20578
rect 6414 20526 6466 20578
rect 7534 20526 7586 20578
rect 7646 20526 7698 20578
rect 13582 20526 13634 20578
rect 17726 20526 17778 20578
rect 17838 20526 17890 20578
rect 17950 20526 18002 20578
rect 18622 20526 18674 20578
rect 21422 20526 21474 20578
rect 23662 20526 23714 20578
rect 28142 20526 28194 20578
rect 28590 20526 28642 20578
rect 29262 20526 29314 20578
rect 30270 20526 30322 20578
rect 32398 20526 32450 20578
rect 32510 20526 32562 20578
rect 32622 20526 32674 20578
rect 36094 20526 36146 20578
rect 39678 20526 39730 20578
rect 39902 20526 39954 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 4734 20190 4786 20242
rect 5742 20190 5794 20242
rect 9662 20190 9714 20242
rect 10334 20190 10386 20242
rect 14030 20190 14082 20242
rect 17726 20190 17778 20242
rect 17838 20190 17890 20242
rect 18622 20190 18674 20242
rect 23438 20190 23490 20242
rect 24446 20190 24498 20242
rect 25230 20190 25282 20242
rect 30606 20190 30658 20242
rect 3614 20078 3666 20130
rect 5182 20078 5234 20130
rect 5630 20078 5682 20130
rect 6414 20078 6466 20130
rect 8206 20078 8258 20130
rect 9774 20078 9826 20130
rect 14142 20078 14194 20130
rect 16718 20078 16770 20130
rect 18062 20078 18114 20130
rect 24222 20078 24274 20130
rect 26238 20078 26290 20130
rect 29150 20078 29202 20130
rect 33406 20078 33458 20130
rect 37662 20078 37714 20130
rect 38446 20078 38498 20130
rect 2718 19966 2770 20018
rect 6190 19966 6242 20018
rect 7310 19966 7362 20018
rect 7870 19966 7922 20018
rect 8430 19966 8482 20018
rect 8654 19966 8706 20018
rect 8878 19966 8930 20018
rect 10446 19966 10498 20018
rect 14702 19966 14754 20018
rect 15038 19966 15090 20018
rect 17390 19966 17442 20018
rect 17614 19966 17666 20018
rect 19854 19966 19906 20018
rect 20526 19966 20578 20018
rect 20974 19966 21026 20018
rect 24782 19966 24834 20018
rect 25566 19966 25618 20018
rect 26574 19966 26626 20018
rect 26686 19966 26738 20018
rect 26798 19966 26850 20018
rect 27246 19966 27298 20018
rect 30382 19966 30434 20018
rect 31950 19966 32002 20018
rect 33630 19966 33682 20018
rect 34078 19966 34130 20018
rect 34974 19966 35026 20018
rect 35310 19966 35362 20018
rect 39006 19966 39058 20018
rect 1934 19854 1986 19906
rect 4062 19854 4114 19906
rect 6526 19854 6578 19906
rect 7086 19854 7138 19906
rect 8766 19854 8818 19906
rect 9550 19854 9602 19906
rect 10894 19854 10946 19906
rect 12238 19854 12290 19906
rect 12686 19854 12738 19906
rect 19182 19854 19234 19906
rect 25790 19854 25842 19906
rect 27582 19854 27634 19906
rect 28030 19854 28082 19906
rect 28478 19854 28530 19906
rect 31502 19854 31554 19906
rect 32510 19854 32562 19906
rect 40014 19854 40066 19906
rect 5854 19742 5906 19794
rect 10334 19742 10386 19794
rect 23998 19742 24050 19794
rect 24558 19742 24610 19794
rect 26126 19742 26178 19794
rect 29710 19742 29762 19794
rect 29934 19742 29986 19794
rect 30158 19742 30210 19794
rect 31054 19742 31106 19794
rect 31278 19742 31330 19794
rect 34414 19742 34466 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 8542 19406 8594 19458
rect 8878 19406 8930 19458
rect 12798 19406 12850 19458
rect 14254 19406 14306 19458
rect 14478 19406 14530 19458
rect 20862 19406 20914 19458
rect 23774 19406 23826 19458
rect 25342 19406 25394 19458
rect 25678 19406 25730 19458
rect 34302 19406 34354 19458
rect 37662 19406 37714 19458
rect 4174 19294 4226 19346
rect 7758 19294 7810 19346
rect 8318 19294 8370 19346
rect 11566 19294 11618 19346
rect 15150 19294 15202 19346
rect 15934 19294 15986 19346
rect 22206 19294 22258 19346
rect 30270 19294 30322 19346
rect 31166 19294 31218 19346
rect 34190 19294 34242 19346
rect 35534 19294 35586 19346
rect 37214 19294 37266 19346
rect 37550 19294 37602 19346
rect 2942 19182 2994 19234
rect 3390 19182 3442 19234
rect 4510 19182 4562 19234
rect 4734 19182 4786 19234
rect 5182 19182 5234 19234
rect 5518 19182 5570 19234
rect 5854 19182 5906 19234
rect 6302 19182 6354 19234
rect 6862 19182 6914 19234
rect 11006 19182 11058 19234
rect 11678 19182 11730 19234
rect 11902 19182 11954 19234
rect 12126 19182 12178 19234
rect 12462 19182 12514 19234
rect 12910 19182 12962 19234
rect 15262 19182 15314 19234
rect 16718 19182 16770 19234
rect 16830 19182 16882 19234
rect 16942 19182 16994 19234
rect 17166 19182 17218 19234
rect 17726 19182 17778 19234
rect 23102 19182 23154 19234
rect 24110 19182 24162 19234
rect 24670 19182 24722 19234
rect 25678 19182 25730 19234
rect 26126 19182 26178 19234
rect 26350 19182 26402 19234
rect 28478 19182 28530 19234
rect 30718 19182 30770 19234
rect 33742 19182 33794 19234
rect 34750 19182 34802 19234
rect 2046 19070 2098 19122
rect 3614 19070 3666 19122
rect 5742 19070 5794 19122
rect 10782 19070 10834 19122
rect 11454 19070 11506 19122
rect 13694 19070 13746 19122
rect 13918 19070 13970 19122
rect 14030 19070 14082 19122
rect 21422 19070 21474 19122
rect 24894 19070 24946 19122
rect 26238 19070 26290 19122
rect 26574 19070 26626 19122
rect 31054 19070 31106 19122
rect 32622 19070 32674 19122
rect 35086 19070 35138 19122
rect 40238 19070 40290 19122
rect 4622 18958 4674 19010
rect 9326 18958 9378 19010
rect 9774 18958 9826 19010
rect 10222 18958 10274 19010
rect 12798 18958 12850 19010
rect 16494 18958 16546 19010
rect 20302 18958 20354 19010
rect 21310 18958 21362 19010
rect 28030 18958 28082 19010
rect 29262 18958 29314 19010
rect 31278 18958 31330 19010
rect 31502 18958 31554 19010
rect 32062 18958 32114 19010
rect 32734 18958 32786 19010
rect 35982 18958 36034 19010
rect 39678 18958 39730 19010
rect 39902 18958 39954 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 4958 18622 5010 18674
rect 5630 18622 5682 18674
rect 6190 18622 6242 18674
rect 7982 18622 8034 18674
rect 8766 18622 8818 18674
rect 13134 18622 13186 18674
rect 13358 18622 13410 18674
rect 15038 18622 15090 18674
rect 15934 18622 15986 18674
rect 17726 18622 17778 18674
rect 18062 18622 18114 18674
rect 18734 18622 18786 18674
rect 24222 18622 24274 18674
rect 24558 18622 24610 18674
rect 6302 18510 6354 18562
rect 6862 18510 6914 18562
rect 6974 18510 7026 18562
rect 7534 18510 7586 18562
rect 8318 18510 8370 18562
rect 12014 18510 12066 18562
rect 14030 18510 14082 18562
rect 14254 18510 14306 18562
rect 14926 18510 14978 18562
rect 15822 18510 15874 18562
rect 22878 18510 22930 18562
rect 2158 18398 2210 18450
rect 2606 18398 2658 18450
rect 8542 18398 8594 18450
rect 8990 18398 9042 18450
rect 9550 18398 9602 18450
rect 10222 18398 10274 18450
rect 10446 18398 10498 18450
rect 11118 18398 11170 18450
rect 13022 18398 13074 18450
rect 13582 18398 13634 18450
rect 15262 18398 15314 18450
rect 15374 18398 15426 18450
rect 16270 18398 16322 18450
rect 17838 18398 17890 18450
rect 18174 18398 18226 18450
rect 19182 18398 19234 18450
rect 19742 18398 19794 18450
rect 21646 18398 21698 18450
rect 23214 18398 23266 18450
rect 23550 18398 23602 18450
rect 25454 18398 25506 18450
rect 26910 18398 26962 18450
rect 33182 18398 33234 18450
rect 33854 18398 33906 18450
rect 8878 18286 8930 18338
rect 12126 18286 12178 18338
rect 12574 18286 12626 18338
rect 13246 18286 13298 18338
rect 13918 18286 13970 18338
rect 16382 18286 16434 18338
rect 16830 18286 16882 18338
rect 20414 18286 20466 18338
rect 21422 18286 21474 18338
rect 21758 18286 21810 18338
rect 21982 18286 22034 18338
rect 22430 18286 22482 18338
rect 23662 18286 23714 18338
rect 25902 18286 25954 18338
rect 26798 18286 26850 18338
rect 27358 18286 27410 18338
rect 27806 18286 27858 18338
rect 28254 18286 28306 18338
rect 28702 18286 28754 18338
rect 29150 18286 29202 18338
rect 29710 18286 29762 18338
rect 30046 18286 30098 18338
rect 30718 18286 30770 18338
rect 31166 18286 31218 18338
rect 31726 18286 31778 18338
rect 32174 18286 32226 18338
rect 34078 18286 34130 18338
rect 34638 18286 34690 18338
rect 35086 18286 35138 18338
rect 35534 18286 35586 18338
rect 6974 18174 7026 18226
rect 11118 18174 11170 18226
rect 11454 18174 11506 18226
rect 11790 18174 11842 18226
rect 12462 18174 12514 18226
rect 23886 18174 23938 18226
rect 24670 18174 24722 18226
rect 28030 18174 28082 18226
rect 28814 18174 28866 18226
rect 31278 18174 31330 18226
rect 32622 18174 32674 18226
rect 34526 18174 34578 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 4958 17838 5010 17890
rect 13470 17838 13522 17890
rect 13806 17838 13858 17890
rect 17502 17838 17554 17890
rect 18174 17838 18226 17890
rect 20414 17838 20466 17890
rect 28030 17838 28082 17890
rect 28254 17838 28306 17890
rect 2270 17726 2322 17778
rect 3166 17726 3218 17778
rect 5070 17726 5122 17778
rect 6190 17726 6242 17778
rect 6526 17726 6578 17778
rect 10670 17726 10722 17778
rect 11454 17726 11506 17778
rect 11902 17726 11954 17778
rect 14142 17726 14194 17778
rect 14254 17726 14306 17778
rect 16270 17726 16322 17778
rect 16606 17726 16658 17778
rect 17054 17726 17106 17778
rect 18062 17726 18114 17778
rect 18398 17726 18450 17778
rect 18958 17726 19010 17778
rect 19966 17726 20018 17778
rect 21870 17726 21922 17778
rect 23214 17726 23266 17778
rect 28030 17726 28082 17778
rect 29374 17726 29426 17778
rect 34638 17726 34690 17778
rect 35982 17726 36034 17778
rect 40014 17726 40066 17778
rect 4734 17614 4786 17666
rect 8878 17614 8930 17666
rect 9550 17614 9602 17666
rect 9774 17614 9826 17666
rect 10782 17614 10834 17666
rect 11790 17614 11842 17666
rect 12126 17614 12178 17666
rect 12238 17614 12290 17666
rect 12574 17614 12626 17666
rect 19854 17614 19906 17666
rect 20302 17614 20354 17666
rect 21310 17614 21362 17666
rect 22766 17614 22818 17666
rect 23998 17614 24050 17666
rect 24670 17614 24722 17666
rect 29710 17614 29762 17666
rect 30382 17614 30434 17666
rect 33854 17614 33906 17666
rect 34302 17614 34354 17666
rect 39118 17614 39170 17666
rect 1710 17502 1762 17554
rect 3726 17502 3778 17554
rect 10110 17502 10162 17554
rect 14366 17502 14418 17554
rect 14926 17502 14978 17554
rect 35534 17502 35586 17554
rect 2606 17390 2658 17442
rect 4062 17390 4114 17442
rect 8542 17390 8594 17442
rect 8990 17390 9042 17442
rect 9102 17390 9154 17442
rect 9998 17390 10050 17442
rect 13582 17390 13634 17442
rect 15374 17390 15426 17442
rect 17502 17390 17554 17442
rect 26910 17390 26962 17442
rect 27694 17390 27746 17442
rect 28478 17390 28530 17442
rect 29486 17390 29538 17442
rect 32846 17390 32898 17442
rect 33406 17390 33458 17442
rect 33630 17390 33682 17442
rect 33742 17390 33794 17442
rect 34526 17390 34578 17442
rect 35086 17390 35138 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 1822 17054 1874 17106
rect 2942 17054 2994 17106
rect 10110 17054 10162 17106
rect 12014 17054 12066 17106
rect 14142 17054 14194 17106
rect 15486 17054 15538 17106
rect 19294 17054 19346 17106
rect 23774 17054 23826 17106
rect 24110 17054 24162 17106
rect 26910 17054 26962 17106
rect 33182 17054 33234 17106
rect 10334 16942 10386 16994
rect 11790 16942 11842 16994
rect 12686 16942 12738 16994
rect 14254 16942 14306 16994
rect 14814 16942 14866 16994
rect 17502 16942 17554 16994
rect 18398 16942 18450 16994
rect 21086 16942 21138 16994
rect 23102 16942 23154 16994
rect 24558 16942 24610 16994
rect 33294 16942 33346 16994
rect 36430 16942 36482 16994
rect 37214 16942 37266 16994
rect 11006 16830 11058 16882
rect 12462 16830 12514 16882
rect 12798 16830 12850 16882
rect 13358 16830 13410 16882
rect 13918 16830 13970 16882
rect 15262 16830 15314 16882
rect 15934 16830 15986 16882
rect 17278 16830 17330 16882
rect 17614 16830 17666 16882
rect 18286 16830 18338 16882
rect 20190 16830 20242 16882
rect 21982 16830 22034 16882
rect 25230 16830 25282 16882
rect 28702 16830 28754 16882
rect 33630 16830 33682 16882
rect 34078 16830 34130 16882
rect 39006 16830 39058 16882
rect 39790 16830 39842 16882
rect 11118 16718 11170 16770
rect 11902 16718 11954 16770
rect 15374 16718 15426 16770
rect 16270 16718 16322 16770
rect 16830 16718 16882 16770
rect 18734 16718 18786 16770
rect 19854 16718 19906 16770
rect 26014 16718 26066 16770
rect 26798 16718 26850 16770
rect 29262 16718 29314 16770
rect 2158 16606 2210 16658
rect 24446 16606 24498 16658
rect 33182 16606 33234 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 10334 16270 10386 16322
rect 12462 16270 12514 16322
rect 12798 16270 12850 16322
rect 13470 16270 13522 16322
rect 18174 16270 18226 16322
rect 34638 16270 34690 16322
rect 36206 16270 36258 16322
rect 12238 16158 12290 16210
rect 13582 16158 13634 16210
rect 14254 16158 14306 16210
rect 19406 16158 19458 16210
rect 20750 16158 20802 16210
rect 26126 16158 26178 16210
rect 31166 16158 31218 16210
rect 32062 16158 32114 16210
rect 35534 16158 35586 16210
rect 36094 16158 36146 16210
rect 2942 16046 2994 16098
rect 6750 16046 6802 16098
rect 7310 16046 7362 16098
rect 14702 16046 14754 16098
rect 15150 16046 15202 16098
rect 19294 16046 19346 16098
rect 21310 16046 21362 16098
rect 21870 16046 21922 16098
rect 25454 16046 25506 16098
rect 28590 16046 28642 16098
rect 29598 16046 29650 16098
rect 31278 16046 31330 16098
rect 31726 16046 31778 16098
rect 32622 16046 32674 16098
rect 32958 16046 33010 16098
rect 33630 16046 33682 16098
rect 34302 16046 34354 16098
rect 39006 16046 39058 16098
rect 2046 15934 2098 15986
rect 12574 15934 12626 15986
rect 19630 15934 19682 15986
rect 25118 15934 25170 15986
rect 27134 15934 27186 15986
rect 27246 15934 27298 15986
rect 28142 15934 28194 15986
rect 29822 15934 29874 15986
rect 30382 15934 30434 15986
rect 31054 15934 31106 15986
rect 33294 15934 33346 15986
rect 33966 15934 34018 15986
rect 34078 15934 34130 15986
rect 34526 15934 34578 15986
rect 40126 15934 40178 15986
rect 9662 15822 9714 15874
rect 10670 15822 10722 15874
rect 17390 15822 17442 15874
rect 24446 15822 24498 15874
rect 26910 15822 26962 15874
rect 27806 15822 27858 15874
rect 29262 15822 29314 15874
rect 32062 15822 32114 15874
rect 32174 15822 32226 15874
rect 32398 15822 32450 15874
rect 33182 15822 33234 15874
rect 33406 15822 33458 15874
rect 35086 15822 35138 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 9662 15486 9714 15538
rect 10110 15486 10162 15538
rect 13582 15486 13634 15538
rect 14142 15486 14194 15538
rect 14366 15486 14418 15538
rect 15598 15486 15650 15538
rect 15822 15486 15874 15538
rect 16830 15486 16882 15538
rect 17502 15486 17554 15538
rect 20078 15486 20130 15538
rect 21758 15486 21810 15538
rect 25790 15486 25842 15538
rect 25902 15486 25954 15538
rect 29486 15486 29538 15538
rect 30270 15486 30322 15538
rect 30718 15486 30770 15538
rect 31614 15486 31666 15538
rect 34638 15486 34690 15538
rect 35534 15486 35586 15538
rect 36094 15486 36146 15538
rect 9550 15374 9602 15426
rect 14478 15374 14530 15426
rect 17614 15374 17666 15426
rect 18510 15374 18562 15426
rect 20862 15374 20914 15426
rect 24110 15374 24162 15426
rect 30494 15374 30546 15426
rect 31950 15374 32002 15426
rect 10670 15262 10722 15314
rect 11118 15262 11170 15314
rect 16270 15262 16322 15314
rect 17278 15262 17330 15314
rect 18734 15262 18786 15314
rect 19182 15262 19234 15314
rect 19406 15262 19458 15314
rect 19630 15262 19682 15314
rect 21758 15262 21810 15314
rect 22094 15262 22146 15314
rect 23326 15262 23378 15314
rect 23774 15262 23826 15314
rect 25678 15262 25730 15314
rect 26350 15262 26402 15314
rect 26686 15262 26738 15314
rect 27246 15262 27298 15314
rect 30942 15262 30994 15314
rect 31054 15262 31106 15314
rect 33294 15262 33346 15314
rect 33630 15262 33682 15314
rect 33854 15262 33906 15314
rect 34078 15262 34130 15314
rect 34414 15262 34466 15314
rect 39006 15262 39058 15314
rect 15374 15150 15426 15202
rect 15710 15150 15762 15202
rect 16718 15150 16770 15202
rect 18062 15150 18114 15202
rect 23214 15150 23266 15202
rect 24446 15150 24498 15202
rect 25230 15150 25282 15202
rect 30830 15150 30882 15202
rect 31502 15150 31554 15202
rect 32510 15150 32562 15202
rect 33406 15150 33458 15202
rect 35086 15150 35138 15202
rect 39790 15150 39842 15202
rect 40350 15150 40402 15202
rect 17950 15038 18002 15090
rect 25342 15038 25394 15090
rect 32062 15038 32114 15090
rect 34750 15038 34802 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 19854 14702 19906 14754
rect 27918 14702 27970 14754
rect 14142 14590 14194 14642
rect 14702 14590 14754 14642
rect 19070 14590 19122 14642
rect 27134 14590 27186 14642
rect 27806 14590 27858 14642
rect 31950 14590 32002 14642
rect 34638 14590 34690 14642
rect 39230 14590 39282 14642
rect 13694 14478 13746 14530
rect 14926 14478 14978 14530
rect 15486 14478 15538 14530
rect 19630 14478 19682 14530
rect 20190 14478 20242 14530
rect 21870 14478 21922 14530
rect 22206 14478 22258 14530
rect 23998 14478 24050 14530
rect 24334 14478 24386 14530
rect 26126 14478 26178 14530
rect 26798 14478 26850 14530
rect 27246 14478 27298 14530
rect 27358 14478 27410 14530
rect 29710 14478 29762 14530
rect 30046 14478 30098 14530
rect 30606 14478 30658 14530
rect 30942 14478 30994 14530
rect 34190 14478 34242 14530
rect 40238 14478 40290 14530
rect 7534 14366 7586 14418
rect 8430 14366 8482 14418
rect 18622 14366 18674 14418
rect 21310 14366 21362 14418
rect 21646 14366 21698 14418
rect 22542 14366 22594 14418
rect 22878 14366 22930 14418
rect 24782 14366 24834 14418
rect 26462 14366 26514 14418
rect 28254 14366 28306 14418
rect 30158 14366 30210 14418
rect 30494 14366 30546 14418
rect 32734 14366 32786 14418
rect 32846 14366 32898 14418
rect 32958 14366 33010 14418
rect 7422 14254 7474 14306
rect 7646 14254 7698 14306
rect 7870 14254 7922 14306
rect 8318 14254 8370 14306
rect 17950 14254 18002 14306
rect 21534 14254 21586 14306
rect 24222 14254 24274 14306
rect 26350 14254 26402 14306
rect 27022 14254 27074 14306
rect 28366 14254 28418 14306
rect 28590 14254 28642 14306
rect 33406 14254 33458 14306
rect 35646 14254 35698 14306
rect 36094 14254 36146 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 16830 13918 16882 13970
rect 19294 13918 19346 13970
rect 21086 13918 21138 13970
rect 24110 13918 24162 13970
rect 26574 13918 26626 13970
rect 33182 13918 33234 13970
rect 38558 13918 38610 13970
rect 5070 13806 5122 13858
rect 8206 13806 8258 13858
rect 13694 13806 13746 13858
rect 16382 13806 16434 13858
rect 17838 13806 17890 13858
rect 19630 13806 19682 13858
rect 20638 13806 20690 13858
rect 22654 13806 22706 13858
rect 27358 13806 27410 13858
rect 28142 13806 28194 13858
rect 30046 13806 30098 13858
rect 30718 13806 30770 13858
rect 32510 13806 32562 13858
rect 33070 13806 33122 13858
rect 33630 13806 33682 13858
rect 37774 13806 37826 13858
rect 5406 13694 5458 13746
rect 8990 13694 9042 13746
rect 15934 13694 15986 13746
rect 19070 13694 19122 13746
rect 20414 13694 20466 13746
rect 21198 13694 21250 13746
rect 21646 13694 21698 13746
rect 22206 13694 22258 13746
rect 25902 13694 25954 13746
rect 26238 13694 26290 13746
rect 26798 13694 26850 13746
rect 27022 13694 27074 13746
rect 27246 13694 27298 13746
rect 27694 13694 27746 13746
rect 28254 13694 28306 13746
rect 28926 13694 28978 13746
rect 30270 13694 30322 13746
rect 31054 13694 31106 13746
rect 31614 13694 31666 13746
rect 32062 13694 32114 13746
rect 32286 13694 32338 13746
rect 33406 13694 33458 13746
rect 34078 13694 34130 13746
rect 34862 13694 34914 13746
rect 35534 13694 35586 13746
rect 39006 13694 39058 13746
rect 6078 13582 6130 13634
rect 9662 13582 9714 13634
rect 21422 13582 21474 13634
rect 23886 13582 23938 13634
rect 25454 13582 25506 13634
rect 27358 13582 27410 13634
rect 27918 13582 27970 13634
rect 31166 13582 31218 13634
rect 32398 13582 32450 13634
rect 34526 13582 34578 13634
rect 40014 13582 40066 13634
rect 21086 13470 21138 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 7198 13134 7250 13186
rect 7310 13134 7362 13186
rect 7534 13134 7586 13186
rect 18846 13134 18898 13186
rect 26014 13134 26066 13186
rect 26910 13134 26962 13186
rect 30158 13134 30210 13186
rect 31278 13134 31330 13186
rect 31838 13134 31890 13186
rect 32510 13134 32562 13186
rect 32734 13134 32786 13186
rect 37774 13134 37826 13186
rect 2942 13022 2994 13074
rect 5070 13022 5122 13074
rect 5630 13022 5682 13074
rect 6526 13022 6578 13074
rect 10894 13022 10946 13074
rect 12014 13022 12066 13074
rect 12462 13022 12514 13074
rect 12910 13022 12962 13074
rect 13694 13022 13746 13074
rect 15262 13022 15314 13074
rect 18510 13022 18562 13074
rect 20414 13022 20466 13074
rect 21646 13022 21698 13074
rect 22878 13022 22930 13074
rect 27134 13022 27186 13074
rect 29262 13022 29314 13074
rect 31502 13022 31554 13074
rect 31950 13022 32002 13074
rect 34190 13022 34242 13074
rect 37326 13022 37378 13074
rect 37662 13022 37714 13074
rect 38670 13022 38722 13074
rect 2270 12910 2322 12962
rect 6078 12910 6130 12962
rect 7982 12910 8034 12962
rect 19070 12910 19122 12962
rect 19406 12910 19458 12962
rect 19742 12910 19794 12962
rect 20638 12910 20690 12962
rect 22094 12910 22146 12962
rect 23662 12910 23714 12962
rect 24782 12910 24834 12962
rect 25230 12910 25282 12962
rect 26686 12910 26738 12962
rect 27806 12910 27858 12962
rect 28030 12910 28082 12962
rect 28366 12910 28418 12962
rect 29150 12910 29202 12962
rect 29822 12910 29874 12962
rect 30046 12910 30098 12962
rect 33070 12910 33122 12962
rect 33182 12910 33234 12962
rect 33406 12910 33458 12962
rect 34078 12910 34130 12962
rect 34750 12910 34802 12962
rect 35310 12910 35362 12962
rect 35758 12910 35810 12962
rect 35982 12910 36034 12962
rect 7646 12798 7698 12850
rect 8766 12798 8818 12850
rect 11230 12798 11282 12850
rect 14366 12798 14418 12850
rect 18286 12798 18338 12850
rect 18510 12798 18562 12850
rect 20414 12798 20466 12850
rect 27582 12798 27634 12850
rect 30830 12798 30882 12850
rect 34974 12798 35026 12850
rect 35646 12798 35698 12850
rect 36318 12798 36370 12850
rect 39454 12798 39506 12850
rect 39678 12798 39730 12850
rect 40238 12798 40290 12850
rect 11342 12686 11394 12738
rect 11454 12686 11506 12738
rect 11902 12686 11954 12738
rect 19630 12686 19682 12738
rect 28142 12686 28194 12738
rect 28254 12686 28306 12738
rect 29374 12686 29426 12738
rect 30158 12686 30210 12738
rect 30942 12686 30994 12738
rect 31166 12686 31218 12738
rect 33294 12686 33346 12738
rect 34302 12686 34354 12738
rect 35086 12686 35138 12738
rect 35422 12686 35474 12738
rect 36206 12686 36258 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4846 12350 4898 12402
rect 18286 12350 18338 12402
rect 20974 12350 21026 12402
rect 27582 12350 27634 12402
rect 30718 12350 30770 12402
rect 32398 12350 32450 12402
rect 34526 12350 34578 12402
rect 8542 12238 8594 12290
rect 14702 12238 14754 12290
rect 18846 12238 18898 12290
rect 19294 12238 19346 12290
rect 21982 12238 22034 12290
rect 22990 12238 23042 12290
rect 25790 12238 25842 12290
rect 28926 12238 28978 12290
rect 30606 12238 30658 12290
rect 31278 12238 31330 12290
rect 33742 12238 33794 12290
rect 34974 12238 35026 12290
rect 5182 12126 5234 12178
rect 13470 12126 13522 12178
rect 13918 12126 13970 12178
rect 17950 12126 18002 12178
rect 19966 12126 20018 12178
rect 20862 12126 20914 12178
rect 22206 12126 22258 12178
rect 23102 12126 23154 12178
rect 25230 12126 25282 12178
rect 28478 12126 28530 12178
rect 29486 12126 29538 12178
rect 30046 12126 30098 12178
rect 30494 12126 30546 12178
rect 33070 12126 33122 12178
rect 33630 12126 33682 12178
rect 34750 12126 34802 12178
rect 5966 12014 6018 12066
rect 8094 12014 8146 12066
rect 10670 12014 10722 12066
rect 12798 12014 12850 12066
rect 16830 12014 16882 12066
rect 18398 12014 18450 12066
rect 20750 12014 20802 12066
rect 22766 12014 22818 12066
rect 27022 12014 27074 12066
rect 28814 12014 28866 12066
rect 34078 12014 34130 12066
rect 34638 12014 34690 12066
rect 35534 12014 35586 12066
rect 35982 12014 36034 12066
rect 17390 11902 17442 11954
rect 17726 11902 17778 11954
rect 18734 11902 18786 11954
rect 19854 11902 19906 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 6862 11566 6914 11618
rect 27246 11566 27298 11618
rect 27806 11566 27858 11618
rect 28254 11566 28306 11618
rect 6974 11454 7026 11506
rect 12910 11454 12962 11506
rect 20526 11454 20578 11506
rect 22654 11454 22706 11506
rect 25342 11454 25394 11506
rect 27358 11454 27410 11506
rect 27694 11454 27746 11506
rect 29710 11454 29762 11506
rect 9438 11342 9490 11394
rect 9998 11342 10050 11394
rect 13582 11342 13634 11394
rect 13918 11342 13970 11394
rect 14926 11342 14978 11394
rect 15598 11342 15650 11394
rect 20414 11342 20466 11394
rect 22878 11342 22930 11394
rect 23774 11342 23826 11394
rect 25454 11342 25506 11394
rect 27918 11342 27970 11394
rect 28478 11342 28530 11394
rect 29598 11342 29650 11394
rect 29934 11342 29986 11394
rect 30046 11342 30098 11394
rect 30494 11342 30546 11394
rect 31166 11342 31218 11394
rect 32062 11342 32114 11394
rect 32846 11342 32898 11394
rect 33406 11342 33458 11394
rect 34190 11342 34242 11394
rect 34526 11342 34578 11394
rect 34750 11342 34802 11394
rect 35646 11342 35698 11394
rect 35870 11342 35922 11394
rect 36206 11342 36258 11394
rect 10782 11230 10834 11282
rect 13470 11230 13522 11282
rect 19406 11230 19458 11282
rect 19742 11230 19794 11282
rect 21870 11230 21922 11282
rect 24446 11230 24498 11282
rect 25118 11230 25170 11282
rect 30942 11230 30994 11282
rect 31054 11230 31106 11282
rect 31278 11230 31330 11282
rect 31726 11230 31778 11282
rect 32734 11230 32786 11282
rect 35086 11230 35138 11282
rect 36094 11230 36146 11282
rect 37214 11230 37266 11282
rect 9662 11118 9714 11170
rect 18062 11118 18114 11170
rect 18622 11118 18674 11170
rect 19070 11118 19122 11170
rect 29262 11118 29314 11170
rect 33966 11118 34018 11170
rect 34302 11118 34354 11170
rect 35198 11118 35250 11170
rect 35310 11118 35362 11170
rect 37774 11118 37826 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 12798 10782 12850 10834
rect 16718 10782 16770 10834
rect 30046 10782 30098 10834
rect 30382 10782 30434 10834
rect 31278 10782 31330 10834
rect 31502 10782 31554 10834
rect 37774 10782 37826 10834
rect 38334 10782 38386 10834
rect 10334 10670 10386 10722
rect 13134 10670 13186 10722
rect 17502 10670 17554 10722
rect 17838 10670 17890 10722
rect 20974 10670 21026 10722
rect 25342 10670 25394 10722
rect 27022 10670 27074 10722
rect 27134 10670 27186 10722
rect 28142 10670 28194 10722
rect 28814 10670 28866 10722
rect 30494 10670 30546 10722
rect 31614 10670 31666 10722
rect 32062 10670 32114 10722
rect 33070 10670 33122 10722
rect 38670 10670 38722 10722
rect 39118 10670 39170 10722
rect 9662 10558 9714 10610
rect 13694 10558 13746 10610
rect 18174 10558 18226 10610
rect 18734 10558 18786 10610
rect 25230 10558 25282 10610
rect 27358 10558 27410 10610
rect 28030 10558 28082 10610
rect 28926 10558 28978 10610
rect 29934 10558 29986 10610
rect 32286 10558 32338 10610
rect 32510 10558 32562 10610
rect 33742 10558 33794 10610
rect 33966 10558 34018 10610
rect 34862 10558 34914 10610
rect 35310 10558 35362 10610
rect 38558 10558 38610 10610
rect 12462 10446 12514 10498
rect 14478 10446 14530 10498
rect 22206 10446 22258 10498
rect 25902 10446 25954 10498
rect 30942 10446 30994 10498
rect 32398 10446 32450 10498
rect 26574 10334 26626 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 10782 9998 10834 10050
rect 11118 9998 11170 10050
rect 14814 9998 14866 10050
rect 19742 9998 19794 10050
rect 29150 9998 29202 10050
rect 29710 9998 29762 10050
rect 29934 9998 29986 10050
rect 34638 9998 34690 10050
rect 11342 9886 11394 9938
rect 12574 9886 12626 9938
rect 13022 9886 13074 9938
rect 13694 9886 13746 9938
rect 13918 9886 13970 9938
rect 15374 9886 15426 9938
rect 19294 9886 19346 9938
rect 19630 9886 19682 9938
rect 20526 9886 20578 9938
rect 21646 9886 21698 9938
rect 22318 9886 22370 9938
rect 20750 9774 20802 9826
rect 21310 9774 21362 9826
rect 22430 9774 22482 9826
rect 24334 9774 24386 9826
rect 24782 9774 24834 9826
rect 25006 9774 25058 9826
rect 26574 9774 26626 9826
rect 30382 9774 30434 9826
rect 30606 9774 30658 9826
rect 32846 9774 32898 9826
rect 14478 9662 14530 9714
rect 20526 9662 20578 9714
rect 23102 9673 23154 9725
rect 26014 9662 26066 9714
rect 27694 9662 27746 9714
rect 28478 9662 28530 9714
rect 28590 9662 28642 9714
rect 29374 9662 29426 9714
rect 32286 9662 32338 9714
rect 33966 9662 34018 9714
rect 34638 9662 34690 9714
rect 14030 9550 14082 9602
rect 14702 9550 14754 9602
rect 24894 9550 24946 9602
rect 25230 9550 25282 9602
rect 27806 9550 27858 9602
rect 28254 9550 28306 9602
rect 30046 9550 30098 9602
rect 30494 9550 30546 9602
rect 30830 9550 30882 9602
rect 34750 9606 34802 9658
rect 31390 9550 31442 9602
rect 33854 9550 33906 9602
rect 35310 9550 35362 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 21310 9214 21362 9266
rect 21870 9214 21922 9266
rect 23214 9214 23266 9266
rect 24782 9214 24834 9266
rect 26798 9214 26850 9266
rect 27358 9214 27410 9266
rect 27582 9214 27634 9266
rect 30382 9214 30434 9266
rect 31950 9214 32002 9266
rect 32174 9214 32226 9266
rect 33406 9214 33458 9266
rect 34078 9214 34130 9266
rect 34638 9214 34690 9266
rect 35086 9214 35138 9266
rect 26014 9102 26066 9154
rect 26462 9102 26514 9154
rect 27022 9102 27074 9154
rect 27134 9102 27186 9154
rect 27694 9102 27746 9154
rect 28590 9102 28642 9154
rect 30270 9102 30322 9154
rect 31502 9102 31554 9154
rect 33854 9102 33906 9154
rect 34190 9102 34242 9154
rect 18174 8990 18226 9042
rect 18846 8990 18898 9042
rect 22430 8990 22482 9042
rect 22654 8990 22706 9042
rect 22878 8990 22930 9042
rect 25678 8990 25730 9042
rect 29150 8990 29202 9042
rect 31614 8990 31666 9042
rect 32062 8990 32114 9042
rect 32622 8990 32674 9042
rect 33070 8990 33122 9042
rect 33406 8990 33458 9042
rect 33742 8990 33794 9042
rect 30942 8878 30994 8930
rect 25342 8766 25394 8818
rect 31502 8766 31554 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 21310 8430 21362 8482
rect 25678 8430 25730 8482
rect 20638 8318 20690 8370
rect 21422 8318 21474 8370
rect 30158 8318 30210 8370
rect 30606 8318 30658 8370
rect 31166 8318 31218 8370
rect 31726 8318 31778 8370
rect 32174 8318 32226 8370
rect 36318 8318 36370 8370
rect 20414 8206 20466 8258
rect 22206 8206 22258 8258
rect 22654 8206 22706 8258
rect 26350 8206 26402 8258
rect 28254 8206 28306 8258
rect 29150 8206 29202 8258
rect 29374 8206 29426 8258
rect 29710 8206 29762 8258
rect 32622 8206 32674 8258
rect 33182 8206 33234 8258
rect 19406 8094 19458 8146
rect 19742 8094 19794 8146
rect 26014 8094 26066 8146
rect 27470 8094 27522 8146
rect 28030 8094 28082 8146
rect 28478 8094 28530 8146
rect 28590 8094 28642 8146
rect 19070 7982 19122 8034
rect 25118 7982 25170 8034
rect 25902 7982 25954 8034
rect 27918 7982 27970 8034
rect 29262 7982 29314 8034
rect 35758 7982 35810 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 21310 7646 21362 7698
rect 22318 7646 22370 7698
rect 26238 7646 26290 7698
rect 26910 7646 26962 7698
rect 27470 7646 27522 7698
rect 27918 7646 27970 7698
rect 33182 7646 33234 7698
rect 35758 7646 35810 7698
rect 23438 7534 23490 7586
rect 23774 7534 23826 7586
rect 28702 7534 28754 7586
rect 31838 7534 31890 7586
rect 31950 7534 32002 7586
rect 32398 7534 32450 7586
rect 35422 7534 35474 7586
rect 35870 7534 35922 7586
rect 18174 7422 18226 7474
rect 18846 7422 18898 7474
rect 30942 7422 30994 7474
rect 31390 7422 31442 7474
rect 25790 7310 25842 7362
rect 25566 7198 25618 7250
rect 26462 7198 26514 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 21310 6862 21362 6914
rect 27470 6862 27522 6914
rect 21422 6750 21474 6802
rect 31838 6750 31890 6802
rect 21982 6638 22034 6690
rect 23774 6638 23826 6690
rect 24446 6638 24498 6690
rect 28366 6638 28418 6690
rect 22430 6414 22482 6466
rect 26798 6414 26850 6466
rect 27918 6414 27970 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 17502 4286 17554 4338
rect 17838 4174 17890 4226
rect 26350 4174 26402 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18846 3614 18898 3666
rect 22206 3614 22258 3666
rect 25678 3614 25730 3666
rect 26910 3614 26962 3666
rect 23102 3502 23154 3554
rect 23550 3502 23602 3554
rect 26126 3502 26178 3554
rect 26462 3502 26514 3554
rect 18398 3390 18450 3442
rect 21758 3390 21810 3442
rect 23326 3390 23378 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 8736 41200 8848 42000
rect 9408 41200 9520 42000
rect 11424 41200 11536 42000
rect 12096 41200 12208 42000
rect 14784 41200 14896 42000
rect 16128 41200 16240 42000
rect 16800 41200 16912 42000
rect 17472 41200 17584 42000
rect 18144 41200 18256 42000
rect 18816 41200 18928 42000
rect 19488 41200 19600 42000
rect 20160 41200 20272 42000
rect 20832 41200 20944 42000
rect 21504 41200 21616 42000
rect 22176 41200 22288 42000
rect 22848 41200 22960 42000
rect 23520 41200 23632 42000
rect 24192 41200 24304 42000
rect 25536 41200 25648 42000
rect 26208 41200 26320 42000
rect 26880 41200 26992 42000
rect 27552 41200 27664 42000
rect 28896 41200 29008 42000
rect 31584 41200 31696 42000
rect 32256 41200 32368 42000
rect 34272 41200 34384 42000
rect 8764 38610 8820 41200
rect 9436 38668 9492 41200
rect 11452 38668 11508 41200
rect 9436 38612 9716 38668
rect 8764 38558 8766 38610
rect 8818 38558 8820 38610
rect 8764 38546 8820 38558
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 9324 37828 9380 37838
rect 8652 37826 9380 37828
rect 8652 37774 9326 37826
rect 9378 37774 9380 37826
rect 8652 37772 9380 37774
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 7532 36484 7588 36494
rect 4060 36372 4116 36382
rect 3948 34130 4004 34142
rect 3948 34078 3950 34130
rect 4002 34078 4004 34130
rect 3948 33908 4004 34078
rect 3948 33842 4004 33852
rect 2044 31668 2100 31678
rect 2044 31574 2100 31612
rect 1708 31556 1764 31566
rect 1708 30996 1764 31500
rect 2492 31556 2548 31566
rect 2492 31462 2548 31500
rect 3276 31556 3332 31566
rect 3276 31218 3332 31500
rect 3276 31166 3278 31218
rect 3330 31166 3332 31218
rect 3276 31154 3332 31166
rect 1708 30930 1764 30940
rect 2828 31108 2884 31118
rect 2492 30772 2548 30782
rect 2828 30772 2884 31052
rect 2492 30770 2884 30772
rect 2492 30718 2494 30770
rect 2546 30718 2884 30770
rect 2492 30716 2884 30718
rect 2492 30706 2548 30716
rect 2156 30212 2212 30222
rect 2156 30118 2212 30156
rect 2828 30210 2884 30716
rect 2828 30158 2830 30210
rect 2882 30158 2884 30210
rect 2828 30146 2884 30158
rect 2044 29538 2100 29550
rect 2044 29486 2046 29538
rect 2098 29486 2100 29538
rect 1708 29426 1764 29438
rect 1708 29374 1710 29426
rect 1762 29374 1764 29426
rect 1708 28980 1764 29374
rect 1708 28914 1764 28924
rect 2044 28868 2100 29486
rect 2492 29314 2548 29326
rect 2492 29262 2494 29314
rect 2546 29262 2548 29314
rect 2492 28980 2548 29262
rect 2492 28914 2548 28924
rect 2044 28802 2100 28812
rect 2940 28756 2996 28766
rect 2940 28642 2996 28700
rect 2940 28590 2942 28642
rect 2994 28590 2996 28642
rect 2940 28578 2996 28590
rect 2156 28420 2212 28430
rect 2156 28326 2212 28364
rect 3836 27860 3892 27870
rect 3836 27766 3892 27804
rect 2828 26290 2884 26302
rect 2828 26238 2830 26290
rect 2882 26238 2884 26290
rect 1932 26178 1988 26190
rect 1932 26126 1934 26178
rect 1986 26126 1988 26178
rect 1932 25620 1988 26126
rect 1932 25554 1988 25564
rect 2156 25282 2212 25294
rect 2156 25230 2158 25282
rect 2210 25230 2212 25282
rect 2044 25060 2100 25070
rect 2044 24946 2100 25004
rect 2044 24894 2046 24946
rect 2098 24894 2100 24946
rect 2044 24882 2100 24894
rect 2156 24948 2212 25230
rect 2156 24882 2212 24892
rect 2828 25284 2884 26238
rect 2940 25620 2996 25630
rect 2940 25506 2996 25564
rect 2940 25454 2942 25506
rect 2994 25454 2996 25506
rect 2940 25442 2996 25454
rect 2828 24946 2884 25228
rect 2828 24894 2830 24946
rect 2882 24894 2884 24946
rect 2828 24882 2884 24894
rect 3612 24948 3668 24958
rect 3612 24854 3668 24892
rect 1708 24722 1764 24734
rect 1708 24670 1710 24722
rect 1762 24670 1764 24722
rect 1708 24276 1764 24670
rect 1708 24210 1764 24220
rect 2492 24610 2548 24622
rect 2492 24558 2494 24610
rect 2546 24558 2548 24610
rect 2492 24276 2548 24558
rect 2492 24210 2548 24220
rect 2268 23940 2324 23950
rect 2268 23846 2324 23884
rect 1708 23714 1764 23726
rect 1708 23662 1710 23714
rect 1762 23662 1764 23714
rect 1708 23604 1764 23662
rect 1708 23538 1764 23548
rect 2716 23714 2772 23726
rect 2716 23662 2718 23714
rect 2770 23662 2772 23714
rect 2716 23604 2772 23662
rect 2716 23538 2772 23548
rect 2828 23380 2884 23390
rect 2828 23154 2884 23324
rect 3388 23380 3444 23390
rect 3388 23286 3444 23324
rect 2828 23102 2830 23154
rect 2882 23102 2884 23154
rect 2828 23090 2884 23102
rect 1932 23044 1988 23054
rect 1932 22950 1988 22988
rect 2828 22370 2884 22382
rect 2828 22318 2830 22370
rect 2882 22318 2884 22370
rect 1932 22260 1988 22270
rect 1932 22166 1988 22204
rect 1596 22148 1652 22158
rect 1596 21810 1652 22092
rect 1596 21758 1598 21810
rect 1650 21758 1652 21810
rect 1596 21746 1652 21758
rect 2156 22146 2212 22158
rect 2156 22094 2158 22146
rect 2210 22094 2212 22146
rect 2156 21588 2212 22094
rect 2828 22148 2884 22318
rect 3836 22370 3892 22382
rect 3836 22318 3838 22370
rect 3890 22318 3892 22370
rect 3276 22260 3332 22270
rect 3276 22166 3332 22204
rect 2828 22082 2884 22092
rect 2380 21812 2436 21822
rect 2380 21718 2436 21756
rect 3836 21700 3892 22318
rect 3836 21634 3892 21644
rect 2156 21522 2212 21532
rect 4060 21588 4116 36316
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 7308 35140 7364 35150
rect 7084 35138 7364 35140
rect 7084 35086 7310 35138
rect 7362 35086 7364 35138
rect 7084 35084 7364 35086
rect 7084 34916 7140 35084
rect 7308 35074 7364 35084
rect 6860 34914 7140 34916
rect 6860 34862 7086 34914
rect 7138 34862 7140 34914
rect 6860 34860 7140 34862
rect 6748 34690 6804 34702
rect 6748 34638 6750 34690
rect 6802 34638 6804 34690
rect 6636 34242 6692 34254
rect 6636 34190 6638 34242
rect 6690 34190 6692 34242
rect 4284 34130 4340 34142
rect 4284 34078 4286 34130
rect 4338 34078 4340 34130
rect 4284 33460 4340 34078
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 6412 33684 6468 33694
rect 4284 33394 4340 33404
rect 6188 33460 6244 33470
rect 6188 33366 6244 33404
rect 6076 33124 6132 33134
rect 6076 33030 6132 33068
rect 6300 33122 6356 33134
rect 6300 33070 6302 33122
rect 6354 33070 6356 33122
rect 6076 32452 6132 32462
rect 5852 32396 6076 32452
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 5852 31890 5908 32396
rect 6076 32358 6132 32396
rect 5852 31838 5854 31890
rect 5906 31838 5908 31890
rect 5852 31826 5908 31838
rect 5964 32116 6020 32126
rect 5740 31556 5796 31566
rect 5740 31462 5796 31500
rect 5628 30994 5684 31006
rect 5628 30942 5630 30994
rect 5682 30942 5684 30994
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5180 29988 5236 29998
rect 5180 29894 5236 29932
rect 5628 29652 5684 30942
rect 5740 29652 5796 29662
rect 5628 29650 5796 29652
rect 5628 29598 5742 29650
rect 5794 29598 5796 29650
rect 5628 29596 5796 29598
rect 5740 29586 5796 29596
rect 5628 29428 5684 29438
rect 5852 29428 5908 29438
rect 5964 29428 6020 32060
rect 6300 32116 6356 33070
rect 6300 32050 6356 32060
rect 6300 31892 6356 31902
rect 6412 31892 6468 33628
rect 6636 33572 6692 34190
rect 6636 33506 6692 33516
rect 6636 33348 6692 33358
rect 6748 33348 6804 34638
rect 6636 33346 6804 33348
rect 6636 33294 6638 33346
rect 6690 33294 6804 33346
rect 6636 33292 6804 33294
rect 6636 33282 6692 33292
rect 6860 32676 6916 34860
rect 7084 34850 7140 34860
rect 7532 35026 7588 36428
rect 7532 34974 7534 35026
rect 7586 34974 7588 35026
rect 6972 34690 7028 34702
rect 6972 34638 6974 34690
rect 7026 34638 7028 34690
rect 6972 34356 7028 34638
rect 7420 34356 7476 34366
rect 6972 34300 7420 34356
rect 7420 34262 7476 34300
rect 7532 33684 7588 34974
rect 7980 35138 8036 35150
rect 7980 35086 7982 35138
rect 8034 35086 8036 35138
rect 7980 35026 8036 35086
rect 8652 35028 8708 37772
rect 9324 37762 9380 37772
rect 9100 37492 9156 37502
rect 9660 37492 9716 38612
rect 9772 38610 9828 38622
rect 11452 38612 11732 38668
rect 9772 38558 9774 38610
rect 9826 38558 9828 38610
rect 9772 38162 9828 38558
rect 9772 38110 9774 38162
rect 9826 38110 9828 38162
rect 9772 38098 9828 38110
rect 11004 38052 11060 38062
rect 11004 37958 11060 37996
rect 11676 38052 11732 38612
rect 12124 38610 12180 41200
rect 12124 38558 12126 38610
rect 12178 38558 12180 38610
rect 12124 38546 12180 38558
rect 13132 38610 13188 38622
rect 13132 38558 13134 38610
rect 13186 38558 13188 38610
rect 12684 38388 12740 38398
rect 12684 38162 12740 38332
rect 13132 38274 13188 38558
rect 13132 38222 13134 38274
rect 13186 38222 13188 38274
rect 13132 38210 13188 38222
rect 14812 38276 14868 41200
rect 15932 38610 15988 38622
rect 15932 38558 15934 38610
rect 15986 38558 15988 38610
rect 14812 38210 14868 38220
rect 15484 38276 15540 38286
rect 15484 38182 15540 38220
rect 12684 38110 12686 38162
rect 12738 38110 12740 38162
rect 12684 38098 12740 38110
rect 11676 37958 11732 37996
rect 11452 37828 11508 37838
rect 11452 37734 11508 37772
rect 12012 37826 12068 37838
rect 12012 37774 12014 37826
rect 12066 37774 12068 37826
rect 9100 37490 9716 37492
rect 9100 37438 9102 37490
rect 9154 37438 9662 37490
rect 9714 37438 9716 37490
rect 9100 37436 9716 37438
rect 9100 37426 9156 37436
rect 9660 37426 9716 37436
rect 11676 37266 11732 37278
rect 11676 37214 11678 37266
rect 11730 37214 11732 37266
rect 10108 37154 10164 37166
rect 10108 37102 10110 37154
rect 10162 37102 10164 37154
rect 9100 36484 9156 36494
rect 9100 36390 9156 36428
rect 9548 36482 9604 36494
rect 9548 36430 9550 36482
rect 9602 36430 9604 36482
rect 9548 35924 9604 36430
rect 9548 35858 9604 35868
rect 7980 34974 7982 35026
rect 8034 34974 8036 35026
rect 7980 34962 8036 34974
rect 8540 35026 8708 35028
rect 8540 34974 8654 35026
rect 8706 34974 8708 35026
rect 8540 34972 8708 34974
rect 8540 34356 8596 34972
rect 8652 34962 8708 34972
rect 9996 35586 10052 35598
rect 9996 35534 9998 35586
rect 10050 35534 10052 35586
rect 8764 34916 8820 34926
rect 8764 34914 9380 34916
rect 8764 34862 8766 34914
rect 8818 34862 9380 34914
rect 8764 34860 9380 34862
rect 8764 34850 8820 34860
rect 9100 34692 9156 34702
rect 7532 33618 7588 33628
rect 8092 34132 8148 34142
rect 6972 33572 7028 33582
rect 6972 33478 7028 33516
rect 8092 33458 8148 34076
rect 8540 34130 8596 34300
rect 8540 34078 8542 34130
rect 8594 34078 8596 34130
rect 8540 34066 8596 34078
rect 8876 34636 9100 34692
rect 8876 34132 8932 34636
rect 9100 34598 9156 34636
rect 9212 34690 9268 34702
rect 9212 34638 9214 34690
rect 9266 34638 9268 34690
rect 8876 34038 8932 34076
rect 9212 34132 9268 34638
rect 9212 34066 9268 34076
rect 9324 34690 9380 34860
rect 9324 34638 9326 34690
rect 9378 34638 9380 34690
rect 8092 33406 8094 33458
rect 8146 33406 8148 33458
rect 8092 33394 8148 33406
rect 8988 34018 9044 34030
rect 8988 33966 8990 34018
rect 9042 33966 9044 34018
rect 7868 33348 7924 33358
rect 7868 33254 7924 33292
rect 8876 33348 8932 33358
rect 8876 33254 8932 33292
rect 7084 33236 7140 33246
rect 7084 33234 7252 33236
rect 7084 33182 7086 33234
rect 7138 33182 7252 33234
rect 7084 33180 7252 33182
rect 7084 33170 7140 33180
rect 6188 31890 6468 31892
rect 6188 31838 6302 31890
rect 6354 31838 6468 31890
rect 6188 31836 6468 31838
rect 6748 32620 6916 32676
rect 6748 31892 6804 32620
rect 6860 32450 6916 32462
rect 6860 32398 6862 32450
rect 6914 32398 6916 32450
rect 6860 32116 6916 32398
rect 6860 32050 6916 32060
rect 7196 32452 7252 33180
rect 8540 33234 8596 33246
rect 8540 33182 8542 33234
rect 8594 33182 8596 33234
rect 8204 33122 8260 33134
rect 8204 33070 8206 33122
rect 8258 33070 8260 33122
rect 8204 32562 8260 33070
rect 8540 32676 8596 33182
rect 8652 33124 8708 33134
rect 8652 33030 8708 33068
rect 8652 32676 8708 32686
rect 8540 32674 8708 32676
rect 8540 32622 8654 32674
rect 8706 32622 8708 32674
rect 8540 32620 8708 32622
rect 8652 32610 8708 32620
rect 8988 32676 9044 33966
rect 9324 33348 9380 34638
rect 9772 34914 9828 34926
rect 9772 34862 9774 34914
rect 9826 34862 9828 34914
rect 9772 33572 9828 34862
rect 9996 34804 10052 35534
rect 9772 33506 9828 33516
rect 9884 34802 10052 34804
rect 9884 34750 9998 34802
rect 10050 34750 10052 34802
rect 9884 34748 10052 34750
rect 9660 33348 9716 33358
rect 9884 33348 9940 34748
rect 9996 34738 10052 34748
rect 10108 34692 10164 37102
rect 10780 37154 10836 37166
rect 10780 37102 10782 37154
rect 10834 37102 10836 37154
rect 10780 36484 10836 37102
rect 11228 37156 11284 37166
rect 11228 37062 11284 37100
rect 10780 36418 10836 36428
rect 11676 36484 11732 37214
rect 12012 36596 12068 37774
rect 13916 37826 13972 37838
rect 13916 37774 13918 37826
rect 13970 37774 13972 37826
rect 12124 37266 12180 37278
rect 12124 37214 12126 37266
rect 12178 37214 12180 37266
rect 12124 36708 12180 37214
rect 12908 37156 12964 37166
rect 12572 36820 12628 36830
rect 12572 36708 12628 36764
rect 12124 36642 12180 36652
rect 12236 36706 12628 36708
rect 12236 36654 12574 36706
rect 12626 36654 12628 36706
rect 12236 36652 12628 36654
rect 11676 36418 11732 36428
rect 11788 36540 12068 36596
rect 11340 35924 11396 35934
rect 11340 35830 11396 35868
rect 11004 35700 11060 35710
rect 11228 35700 11284 35710
rect 11004 35606 11060 35644
rect 11116 35698 11284 35700
rect 11116 35646 11230 35698
rect 11282 35646 11284 35698
rect 11116 35644 11284 35646
rect 10556 35588 10612 35598
rect 10444 35586 10612 35588
rect 10444 35534 10558 35586
rect 10610 35534 10612 35586
rect 10444 35532 10612 35534
rect 10108 34468 10164 34636
rect 9996 34412 10164 34468
rect 10220 34690 10276 34702
rect 10220 34638 10222 34690
rect 10274 34638 10276 34690
rect 9996 33458 10052 34412
rect 10108 34132 10164 34142
rect 10108 34038 10164 34076
rect 10220 33906 10276 34638
rect 10444 34690 10500 35532
rect 10556 35522 10612 35532
rect 11116 35140 11172 35644
rect 11228 35634 11284 35644
rect 11452 35700 11508 35710
rect 11452 35606 11508 35644
rect 10556 35084 11172 35140
rect 11676 35252 11732 35262
rect 10556 35026 10612 35084
rect 10556 34974 10558 35026
rect 10610 34974 10612 35026
rect 10556 34962 10612 34974
rect 10892 34972 11396 35028
rect 10668 34916 10724 34926
rect 10892 34916 10948 34972
rect 10668 34914 10948 34916
rect 10668 34862 10670 34914
rect 10722 34862 10948 34914
rect 10668 34860 10948 34862
rect 10668 34850 10724 34860
rect 10444 34638 10446 34690
rect 10498 34638 10500 34690
rect 10220 33854 10222 33906
rect 10274 33854 10276 33906
rect 10220 33842 10276 33854
rect 10332 34020 10388 34030
rect 9996 33406 9998 33458
rect 10050 33406 10052 33458
rect 9996 33394 10052 33406
rect 9324 33346 9716 33348
rect 9324 33294 9662 33346
rect 9714 33294 9716 33346
rect 9324 33292 9716 33294
rect 9660 33282 9716 33292
rect 9772 33292 9940 33348
rect 10108 33348 10164 33358
rect 10164 33292 10276 33348
rect 9100 33234 9156 33246
rect 9100 33182 9102 33234
rect 9154 33182 9156 33234
rect 9100 32788 9156 33182
rect 9100 32722 9156 32732
rect 9548 33122 9604 33134
rect 9548 33070 9550 33122
rect 9602 33070 9604 33122
rect 8988 32610 9044 32620
rect 8204 32510 8206 32562
rect 8258 32510 8260 32562
rect 7308 32452 7364 32462
rect 7252 32450 7364 32452
rect 7252 32398 7310 32450
rect 7362 32398 7364 32450
rect 7252 32396 7364 32398
rect 6860 31892 6916 31902
rect 6748 31890 6916 31892
rect 6748 31838 6862 31890
rect 6914 31838 6916 31890
rect 6748 31836 6916 31838
rect 6188 30994 6244 31836
rect 6300 31826 6356 31836
rect 6524 31108 6580 31118
rect 6524 31014 6580 31052
rect 6636 31108 6692 31118
rect 6748 31108 6804 31836
rect 6860 31826 6916 31836
rect 7196 31444 7252 32396
rect 7308 32386 7364 32396
rect 7756 32450 7812 32462
rect 7756 32398 7758 32450
rect 7810 32398 7812 32450
rect 7756 32002 7812 32398
rect 7756 31950 7758 32002
rect 7810 31950 7812 32002
rect 7756 31938 7812 31950
rect 8204 31892 8260 32510
rect 8204 31826 8260 31836
rect 7756 31778 7812 31790
rect 7756 31726 7758 31778
rect 7810 31726 7812 31778
rect 7308 31668 7364 31678
rect 7308 31574 7364 31612
rect 7756 31668 7812 31726
rect 9548 31780 9604 33070
rect 9548 31714 9604 31724
rect 7420 31554 7476 31566
rect 7420 31502 7422 31554
rect 7474 31502 7476 31554
rect 7196 31388 7364 31444
rect 6636 31106 6916 31108
rect 6636 31054 6638 31106
rect 6690 31054 6916 31106
rect 6636 31052 6916 31054
rect 6636 31042 6692 31052
rect 6188 30942 6190 30994
rect 6242 30942 6244 30994
rect 6076 30212 6132 30222
rect 6076 30118 6132 30156
rect 6188 29652 6244 30942
rect 6524 30772 6580 30782
rect 6412 30770 6580 30772
rect 6412 30718 6526 30770
rect 6578 30718 6580 30770
rect 6412 30716 6580 30718
rect 6300 30098 6356 30110
rect 6300 30046 6302 30098
rect 6354 30046 6356 30098
rect 6300 29988 6356 30046
rect 6300 29922 6356 29932
rect 6188 29596 6356 29652
rect 5628 29334 5684 29372
rect 5740 29426 6132 29428
rect 5740 29374 5854 29426
rect 5906 29374 6132 29426
rect 5740 29372 6132 29374
rect 5292 29314 5348 29326
rect 5292 29262 5294 29314
rect 5346 29262 5348 29314
rect 5292 29204 5348 29262
rect 5740 29204 5796 29372
rect 5852 29362 5908 29372
rect 5292 29148 5796 29204
rect 6076 29316 6132 29372
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4284 28420 4340 28430
rect 4284 27858 4340 28364
rect 5852 28418 5908 28430
rect 5852 28366 5854 28418
rect 5906 28366 5908 28418
rect 5852 28196 5908 28366
rect 5964 28420 6020 28430
rect 5964 28326 6020 28364
rect 6076 28418 6132 29260
rect 6188 29426 6244 29438
rect 6188 29374 6190 29426
rect 6242 29374 6244 29426
rect 6188 29314 6244 29374
rect 6188 29262 6190 29314
rect 6242 29262 6244 29314
rect 6188 29250 6244 29262
rect 6300 28644 6356 29596
rect 6412 29314 6468 30716
rect 6524 30706 6580 30716
rect 6748 30212 6804 30222
rect 6748 30118 6804 30156
rect 6524 30100 6580 30110
rect 6524 30006 6580 30044
rect 6636 29986 6692 29998
rect 6636 29934 6638 29986
rect 6690 29934 6692 29986
rect 6636 29540 6692 29934
rect 6860 29652 6916 31052
rect 7196 30884 7252 30894
rect 6972 30882 7252 30884
rect 6972 30830 7198 30882
rect 7250 30830 7252 30882
rect 6972 30828 7252 30830
rect 6972 30210 7028 30828
rect 7196 30818 7252 30828
rect 7308 30324 7364 31388
rect 7420 31108 7476 31502
rect 7420 31042 7476 31052
rect 7756 30996 7812 31612
rect 8092 31666 8148 31678
rect 8092 31614 8094 31666
rect 8146 31614 8148 31666
rect 8092 31556 8148 31614
rect 8876 31668 8932 31678
rect 8932 31612 9044 31668
rect 8876 31574 8932 31612
rect 8540 31556 8596 31566
rect 8092 31554 8596 31556
rect 8092 31502 8542 31554
rect 8594 31502 8596 31554
rect 8092 31500 8596 31502
rect 7532 30994 7812 30996
rect 7532 30942 7758 30994
rect 7810 30942 7812 30994
rect 7532 30940 7812 30942
rect 7308 30268 7476 30324
rect 6972 30158 6974 30210
rect 7026 30158 7028 30210
rect 6972 30146 7028 30158
rect 7308 30100 7364 30110
rect 7308 30006 7364 30044
rect 7084 29652 7140 29662
rect 6860 29650 7140 29652
rect 6860 29598 7086 29650
rect 7138 29598 7140 29650
rect 6860 29596 7140 29598
rect 6636 29474 6692 29484
rect 6412 29262 6414 29314
rect 6466 29262 6468 29314
rect 6412 29250 6468 29262
rect 6636 29316 6692 29326
rect 6636 29222 6692 29260
rect 6860 28756 6916 28766
rect 6076 28366 6078 28418
rect 6130 28366 6132 28418
rect 5852 28130 5908 28140
rect 4284 27806 4286 27858
rect 4338 27806 4340 27858
rect 4284 27794 4340 27806
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 6076 26908 6132 28366
rect 6188 28588 6356 28644
rect 6412 28644 6468 28654
rect 6636 28644 6692 28654
rect 6412 28642 6692 28644
rect 6412 28590 6414 28642
rect 6466 28590 6638 28642
rect 6690 28590 6692 28642
rect 6412 28588 6692 28590
rect 6188 27860 6244 28588
rect 6412 28578 6468 28588
rect 6636 28578 6692 28588
rect 6860 28530 6916 28700
rect 6860 28478 6862 28530
rect 6914 28478 6916 28530
rect 6860 28466 6916 28478
rect 6972 28642 7028 29596
rect 7084 29586 7140 29596
rect 6972 28590 6974 28642
rect 7026 28590 7028 28642
rect 6748 28084 6804 28094
rect 6748 27990 6804 28028
rect 6188 27794 6244 27804
rect 6300 26964 6356 26974
rect 5852 26852 6356 26908
rect 5628 26180 5684 26190
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4732 25508 4788 25518
rect 5068 25508 5124 25518
rect 4732 25506 5124 25508
rect 4732 25454 4734 25506
rect 4786 25454 5070 25506
rect 5122 25454 5124 25506
rect 4732 25452 5124 25454
rect 4732 25442 4788 25452
rect 4956 25282 5012 25294
rect 4956 25230 4958 25282
rect 5010 25230 5012 25282
rect 4956 24948 5012 25230
rect 4956 24882 5012 24892
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4844 22484 4900 22494
rect 5068 22484 5124 25452
rect 5628 25506 5684 26124
rect 5628 25454 5630 25506
rect 5682 25454 5684 25506
rect 5628 25442 5684 25454
rect 5852 25508 5908 26852
rect 6300 26516 6356 26852
rect 6412 26516 6468 26526
rect 6300 26514 6468 26516
rect 6300 26462 6414 26514
rect 6466 26462 6468 26514
rect 6300 26460 6468 26462
rect 6412 26450 6468 26460
rect 6972 26178 7028 28590
rect 7308 28756 7364 28766
rect 7308 28082 7364 28700
rect 7308 28030 7310 28082
rect 7362 28030 7364 28082
rect 7308 28018 7364 28030
rect 6972 26126 6974 26178
rect 7026 26126 7028 26178
rect 6748 25844 6804 25854
rect 6972 25844 7028 26126
rect 6804 25788 7028 25844
rect 7084 27860 7140 27870
rect 7084 27188 7140 27804
rect 7420 27748 7476 30268
rect 7532 29426 7588 30940
rect 7756 30930 7812 30940
rect 7980 30996 8036 31006
rect 7532 29374 7534 29426
rect 7586 29374 7588 29426
rect 7532 29362 7588 29374
rect 7644 29540 7700 29550
rect 7644 28756 7700 29484
rect 7980 29426 8036 30940
rect 8092 30994 8148 31500
rect 8540 31490 8596 31500
rect 8764 31554 8820 31566
rect 8764 31502 8766 31554
rect 8818 31502 8820 31554
rect 8764 31332 8820 31502
rect 8092 30942 8094 30994
rect 8146 30942 8148 30994
rect 8092 30930 8148 30942
rect 8428 31276 8764 31332
rect 8092 30322 8148 30334
rect 8092 30270 8094 30322
rect 8146 30270 8148 30322
rect 8092 29764 8148 30270
rect 8204 30212 8260 30222
rect 8316 30212 8372 30222
rect 8204 30210 8316 30212
rect 8204 30158 8206 30210
rect 8258 30158 8316 30210
rect 8204 30156 8316 30158
rect 8428 30212 8484 31276
rect 8764 31266 8820 31276
rect 8540 31108 8596 31118
rect 8764 31108 8820 31118
rect 8540 31014 8596 31052
rect 8652 31106 8820 31108
rect 8652 31054 8766 31106
rect 8818 31054 8820 31106
rect 8652 31052 8820 31054
rect 8652 30996 8708 31052
rect 8764 31042 8820 31052
rect 8652 30930 8708 30940
rect 8876 30882 8932 30894
rect 8876 30830 8878 30882
rect 8930 30830 8932 30882
rect 8428 30156 8820 30212
rect 8204 30146 8260 30156
rect 8092 29698 8148 29708
rect 8316 29540 8372 30156
rect 8540 29988 8596 29998
rect 8428 29540 8484 29550
rect 8316 29538 8484 29540
rect 8316 29486 8430 29538
rect 8482 29486 8484 29538
rect 8316 29484 8484 29486
rect 8428 29474 8484 29484
rect 7980 29374 7982 29426
rect 8034 29374 8036 29426
rect 7980 29362 8036 29374
rect 7644 28642 7700 28700
rect 8316 28756 8372 28766
rect 8316 28662 8372 28700
rect 7644 28590 7646 28642
rect 7698 28590 7700 28642
rect 7644 28578 7700 28590
rect 8204 28644 8260 28654
rect 8204 28550 8260 28588
rect 7532 28084 7588 28094
rect 7532 27990 7588 28028
rect 7644 27748 7700 27758
rect 8092 27748 8148 27758
rect 7420 27746 8148 27748
rect 7420 27694 7646 27746
rect 7698 27694 8094 27746
rect 8146 27694 8148 27746
rect 7420 27692 8148 27694
rect 7644 27682 7700 27692
rect 8092 27636 8148 27692
rect 8092 27570 8148 27580
rect 7420 27188 7476 27198
rect 7084 27186 7476 27188
rect 7084 27134 7422 27186
rect 7474 27134 7476 27186
rect 7084 27132 7476 27134
rect 6188 25508 6244 25518
rect 6412 25508 6468 25518
rect 5852 25506 6020 25508
rect 5852 25454 5854 25506
rect 5906 25454 6020 25506
rect 5852 25452 6020 25454
rect 5852 25442 5908 25452
rect 5740 25282 5796 25294
rect 5740 25230 5742 25282
rect 5794 25230 5796 25282
rect 5404 24724 5460 24734
rect 5740 24724 5796 25230
rect 5852 24724 5908 24734
rect 5740 24722 5908 24724
rect 5740 24670 5854 24722
rect 5906 24670 5908 24722
rect 5740 24668 5908 24670
rect 5404 23380 5460 24668
rect 5852 24658 5908 24668
rect 4844 22482 5068 22484
rect 4844 22430 4846 22482
rect 4898 22430 5068 22482
rect 4844 22428 5068 22430
rect 4844 22418 4900 22428
rect 4732 22146 4788 22158
rect 4732 22094 4734 22146
rect 4786 22094 4788 22146
rect 4732 21812 4788 22094
rect 4732 21746 4788 21756
rect 4060 21522 4116 21532
rect 4732 21588 4788 21598
rect 4732 21586 4900 21588
rect 4732 21534 4734 21586
rect 4786 21534 4900 21586
rect 4732 21532 4900 21534
rect 4732 21522 4788 21532
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4508 21028 4564 21038
rect 1708 20916 1764 20926
rect 1708 20802 1764 20860
rect 3724 20916 3780 20926
rect 3724 20822 3780 20860
rect 1708 20750 1710 20802
rect 1762 20750 1764 20802
rect 1708 20738 1764 20750
rect 4284 20804 4340 20814
rect 4284 20710 4340 20748
rect 4508 20802 4564 20972
rect 4620 20916 4676 20926
rect 4844 20916 4900 21532
rect 4620 20914 4900 20916
rect 4620 20862 4622 20914
rect 4674 20862 4900 20914
rect 4620 20860 4900 20862
rect 4620 20850 4676 20860
rect 4508 20750 4510 20802
rect 4562 20750 4564 20802
rect 4508 20738 4564 20750
rect 2268 20690 2324 20702
rect 2268 20638 2270 20690
rect 2322 20638 2324 20690
rect 2268 20132 2324 20638
rect 3164 20690 3220 20702
rect 3164 20638 3166 20690
rect 3218 20638 3220 20690
rect 2604 20578 2660 20590
rect 2604 20526 2606 20578
rect 2658 20526 2660 20578
rect 2604 20244 2660 20526
rect 2604 20178 2660 20188
rect 2268 20066 2324 20076
rect 2716 20018 2772 20030
rect 2716 19966 2718 20018
rect 2770 19966 2772 20018
rect 1932 19906 1988 19918
rect 1932 19854 1934 19906
rect 1986 19854 1988 19906
rect 1932 19572 1988 19854
rect 1932 19506 1988 19516
rect 2044 19124 2100 19134
rect 2044 19030 2100 19068
rect 2716 18564 2772 19966
rect 3164 19796 3220 20638
rect 4732 20692 4788 20702
rect 3612 20244 3668 20254
rect 3612 20130 3668 20188
rect 4732 20244 4788 20636
rect 4732 20242 4900 20244
rect 4732 20190 4734 20242
rect 4786 20190 4900 20242
rect 4732 20188 4900 20190
rect 4732 20178 4788 20188
rect 3612 20078 3614 20130
rect 3666 20078 3668 20130
rect 3612 20066 3668 20078
rect 4172 20132 4228 20142
rect 4060 19908 4116 19918
rect 3164 19730 3220 19740
rect 3388 19906 4116 19908
rect 3388 19854 4062 19906
rect 4114 19854 4116 19906
rect 3388 19852 4116 19854
rect 2940 19236 2996 19246
rect 2940 19142 2996 19180
rect 3388 19234 3444 19852
rect 4060 19842 4116 19852
rect 3388 19182 3390 19234
rect 3442 19182 3444 19234
rect 2716 18498 2772 18508
rect 3164 19012 3220 19022
rect 2156 18452 2212 18462
rect 1708 17556 1764 17566
rect 1764 17500 1876 17556
rect 1708 17462 1764 17500
rect 1820 17106 1876 17500
rect 1820 17054 1822 17106
rect 1874 17054 1876 17106
rect 1820 17042 1876 17054
rect 2156 16884 2212 18396
rect 2604 18450 2660 18462
rect 2604 18398 2606 18450
rect 2658 18398 2660 18450
rect 2604 18340 2660 18398
rect 2604 18274 2660 18284
rect 2268 18228 2324 18238
rect 2268 17778 2324 18172
rect 2268 17726 2270 17778
rect 2322 17726 2324 17778
rect 2268 17714 2324 17726
rect 3164 17778 3220 18956
rect 3388 18116 3444 19182
rect 4172 19346 4228 20076
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4172 19294 4174 19346
rect 4226 19294 4228 19346
rect 3612 19124 3668 19134
rect 3612 19030 3668 19068
rect 4172 19012 4228 19294
rect 4508 19348 4564 19358
rect 4508 19234 4564 19292
rect 4508 19182 4510 19234
rect 4562 19182 4564 19234
rect 4508 19170 4564 19182
rect 4732 19236 4788 19246
rect 4844 19236 4900 20188
rect 4732 19234 4900 19236
rect 4732 19182 4734 19234
rect 4786 19182 4900 19234
rect 4732 19180 4900 19182
rect 4732 19170 4788 19180
rect 4172 18946 4228 18956
rect 4620 19010 4676 19022
rect 4620 18958 4622 19010
rect 4674 18958 4676 19010
rect 3388 18050 3444 18060
rect 3724 18564 3780 18574
rect 3164 17726 3166 17778
rect 3218 17726 3220 17778
rect 3164 17714 3220 17726
rect 3724 17556 3780 18508
rect 4620 18340 4676 18958
rect 4620 18274 4676 18284
rect 4956 18674 5012 18686
rect 4956 18622 4958 18674
rect 5010 18622 5012 18674
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4956 17890 5012 18622
rect 4956 17838 4958 17890
rect 5010 17838 5012 17890
rect 4956 17826 5012 17838
rect 5068 17778 5124 22428
rect 5292 23378 5460 23380
rect 5292 23326 5406 23378
rect 5458 23326 5460 23378
rect 5292 23324 5460 23326
rect 5292 21586 5348 23324
rect 5404 23314 5460 23324
rect 5740 22484 5796 22494
rect 5740 22390 5796 22428
rect 5628 22148 5684 22158
rect 5628 21810 5684 22092
rect 5628 21758 5630 21810
rect 5682 21758 5684 21810
rect 5628 21746 5684 21758
rect 5740 21812 5796 21822
rect 5740 21698 5796 21756
rect 5740 21646 5742 21698
rect 5794 21646 5796 21698
rect 5292 21534 5294 21586
rect 5346 21534 5348 21586
rect 5292 21522 5348 21534
rect 5404 21586 5460 21598
rect 5404 21534 5406 21586
rect 5458 21534 5460 21586
rect 5180 20804 5236 20814
rect 5404 20804 5460 21534
rect 5180 20802 5460 20804
rect 5180 20750 5182 20802
rect 5234 20750 5460 20802
rect 5180 20748 5460 20750
rect 5180 20738 5236 20748
rect 5740 20580 5796 21646
rect 5964 20804 6020 25452
rect 6188 25506 6468 25508
rect 6188 25454 6190 25506
rect 6242 25454 6414 25506
rect 6466 25454 6468 25506
rect 6188 25452 6468 25454
rect 6188 25442 6244 25452
rect 6412 25442 6468 25452
rect 6748 25506 6804 25788
rect 6748 25454 6750 25506
rect 6802 25454 6804 25506
rect 6636 25284 6692 25294
rect 6636 25190 6692 25228
rect 6524 24724 6580 24734
rect 6524 24630 6580 24668
rect 6748 22482 6804 25454
rect 6860 24948 6916 24958
rect 7084 24948 7140 27132
rect 7420 27122 7476 27132
rect 8540 27188 8596 29932
rect 8764 29538 8820 30156
rect 8876 30210 8932 30830
rect 8876 30158 8878 30210
rect 8930 30158 8932 30210
rect 8876 30146 8932 30158
rect 8764 29486 8766 29538
rect 8818 29486 8820 29538
rect 8652 28868 8708 28878
rect 8652 27970 8708 28812
rect 8764 28644 8820 29486
rect 8876 29540 8932 29550
rect 8876 29446 8932 29484
rect 8988 28980 9044 31612
rect 9212 31666 9268 31678
rect 9212 31614 9214 31666
rect 9266 31614 9268 31666
rect 9212 31108 9268 31614
rect 9212 31042 9268 31052
rect 9324 31554 9380 31566
rect 9548 31556 9604 31566
rect 9324 31502 9326 31554
rect 9378 31502 9380 31554
rect 9324 30996 9380 31502
rect 9324 30930 9380 30940
rect 9436 31554 9604 31556
rect 9436 31502 9550 31554
rect 9602 31502 9604 31554
rect 9436 31500 9604 31502
rect 9324 30210 9380 30222
rect 9324 30158 9326 30210
rect 9378 30158 9380 30210
rect 9100 29652 9156 29662
rect 9324 29652 9380 30158
rect 9436 30098 9492 31500
rect 9548 31490 9604 31500
rect 9548 31332 9604 31342
rect 9548 31106 9604 31276
rect 9548 31054 9550 31106
rect 9602 31054 9604 31106
rect 9548 31042 9604 31054
rect 9660 31108 9716 31118
rect 9660 30994 9716 31052
rect 9660 30942 9662 30994
rect 9714 30942 9716 30994
rect 9660 30930 9716 30942
rect 9772 30772 9828 33292
rect 10108 33282 10164 33292
rect 10108 33124 10164 33134
rect 9884 32788 9940 32798
rect 9940 32732 10052 32788
rect 9884 32722 9940 32732
rect 9996 32674 10052 32732
rect 9996 32622 9998 32674
rect 10050 32622 10052 32674
rect 9996 32610 10052 32622
rect 10108 32676 10164 33068
rect 9884 32564 9940 32574
rect 9884 32470 9940 32508
rect 10108 32562 10164 32620
rect 10108 32510 10110 32562
rect 10162 32510 10164 32562
rect 10108 32498 10164 32510
rect 9884 31892 9940 31902
rect 9884 30994 9940 31836
rect 9884 30942 9886 30994
rect 9938 30942 9940 30994
rect 9884 30930 9940 30942
rect 10108 31668 10164 31678
rect 10108 30994 10164 31612
rect 10108 30942 10110 30994
rect 10162 30942 10164 30994
rect 10108 30930 10164 30942
rect 9436 30046 9438 30098
rect 9490 30046 9492 30098
rect 9436 30034 9492 30046
rect 9548 30716 9828 30772
rect 9548 29988 9604 30716
rect 10220 30436 10276 33292
rect 10332 31220 10388 33964
rect 10444 33908 10500 34638
rect 11004 34802 11060 34814
rect 11004 34750 11006 34802
rect 11058 34750 11060 34802
rect 10780 34130 10836 34142
rect 10780 34078 10782 34130
rect 10834 34078 10836 34130
rect 10780 34020 10836 34078
rect 11004 34020 11060 34750
rect 11340 34242 11396 34972
rect 11676 34914 11732 35196
rect 11676 34862 11678 34914
rect 11730 34862 11732 34914
rect 11676 34850 11732 34862
rect 11788 34916 11844 36540
rect 11900 36260 11956 36270
rect 11900 36166 11956 36204
rect 12236 35922 12292 36652
rect 12572 36642 12628 36652
rect 12908 36596 12964 37100
rect 13916 36820 13972 37774
rect 14812 37826 14868 37838
rect 14812 37774 14814 37826
rect 14866 37774 14868 37826
rect 14588 37492 14644 37502
rect 14588 37490 14756 37492
rect 14588 37438 14590 37490
rect 14642 37438 14756 37490
rect 14588 37436 14756 37438
rect 14588 37426 14644 37436
rect 13916 36754 13972 36764
rect 12908 36502 12964 36540
rect 13468 36708 13524 36718
rect 13132 36484 13188 36494
rect 12796 36260 12852 36270
rect 12796 36166 12852 36204
rect 13132 35924 13188 36428
rect 13468 36370 13524 36652
rect 13468 36318 13470 36370
rect 13522 36318 13524 36370
rect 13468 36306 13524 36318
rect 13580 36596 13636 36606
rect 12236 35870 12238 35922
rect 12290 35870 12292 35922
rect 12012 35810 12068 35822
rect 12012 35758 12014 35810
rect 12066 35758 12068 35810
rect 11900 35700 11956 35710
rect 12012 35700 12068 35758
rect 11900 35698 12068 35700
rect 11900 35646 11902 35698
rect 11954 35646 12068 35698
rect 11900 35644 12068 35646
rect 11900 35634 11956 35644
rect 12236 35364 12292 35870
rect 12908 35922 13188 35924
rect 12908 35870 13134 35922
rect 13186 35870 13188 35922
rect 12908 35868 13188 35870
rect 11900 34916 11956 34926
rect 11788 34914 11956 34916
rect 11788 34862 11902 34914
rect 11954 34862 11956 34914
rect 11788 34860 11956 34862
rect 11340 34190 11342 34242
rect 11394 34190 11396 34242
rect 11340 34178 11396 34190
rect 11452 34130 11508 34142
rect 11452 34078 11454 34130
rect 11506 34078 11508 34130
rect 11452 34020 11508 34078
rect 11900 34132 11956 34860
rect 11900 34066 11956 34076
rect 12012 34130 12068 34142
rect 12012 34078 12014 34130
rect 12066 34078 12068 34130
rect 10780 33964 11396 34020
rect 10444 33852 11284 33908
rect 10556 33572 10612 33582
rect 10612 33516 10724 33572
rect 10556 33478 10612 33516
rect 10668 32788 10724 33516
rect 10892 33346 10948 33358
rect 10892 33294 10894 33346
rect 10946 33294 10948 33346
rect 10892 32900 10948 33294
rect 11116 33234 11172 33246
rect 11116 33182 11118 33234
rect 11170 33182 11172 33234
rect 11116 33124 11172 33182
rect 11116 33058 11172 33068
rect 10892 32844 11172 32900
rect 10668 32732 10836 32788
rect 10444 32676 10500 32686
rect 10444 32674 10724 32676
rect 10444 32622 10446 32674
rect 10498 32622 10724 32674
rect 10444 32620 10724 32622
rect 10444 32610 10500 32620
rect 10668 32562 10724 32620
rect 10668 32510 10670 32562
rect 10722 32510 10724 32562
rect 10668 32498 10724 32510
rect 10780 32452 10836 32732
rect 10892 32676 10948 32686
rect 10892 32582 10948 32620
rect 11004 32562 11060 32574
rect 11004 32510 11006 32562
rect 11058 32510 11060 32562
rect 11004 32452 11060 32510
rect 10780 32396 11060 32452
rect 11116 32564 11172 32844
rect 10556 31220 10612 31230
rect 10332 31218 10612 31220
rect 10332 31166 10558 31218
rect 10610 31166 10612 31218
rect 10332 31164 10612 31166
rect 10556 31154 10612 31164
rect 11116 31218 11172 32508
rect 11116 31166 11118 31218
rect 11170 31166 11172 31218
rect 11116 31154 11172 31166
rect 11004 30994 11060 31006
rect 11004 30942 11006 30994
rect 11058 30942 11060 30994
rect 10220 30380 10388 30436
rect 9772 30324 9828 30334
rect 9772 30230 9828 30268
rect 10220 30212 10276 30222
rect 10220 30118 10276 30156
rect 9548 29922 9604 29932
rect 9100 29650 9324 29652
rect 9100 29598 9102 29650
rect 9154 29598 9324 29650
rect 9100 29596 9324 29598
rect 9100 29586 9156 29596
rect 9324 29558 9380 29596
rect 10220 29764 10276 29774
rect 10220 29650 10276 29708
rect 10220 29598 10222 29650
rect 10274 29598 10276 29650
rect 10220 29586 10276 29598
rect 9884 29538 9940 29550
rect 9884 29486 9886 29538
rect 9938 29486 9940 29538
rect 9772 29426 9828 29438
rect 9772 29374 9774 29426
rect 9826 29374 9828 29426
rect 8988 28924 9268 28980
rect 9212 28754 9268 28924
rect 9212 28702 9214 28754
rect 9266 28702 9268 28754
rect 8988 28644 9044 28654
rect 8820 28642 9044 28644
rect 8820 28590 8990 28642
rect 9042 28590 9044 28642
rect 8820 28588 9044 28590
rect 8764 28082 8820 28588
rect 8988 28578 9044 28588
rect 8764 28030 8766 28082
rect 8818 28030 8820 28082
rect 8764 28018 8820 28030
rect 8652 27918 8654 27970
rect 8706 27918 8708 27970
rect 8652 27906 8708 27918
rect 9212 27300 9268 28702
rect 9772 28756 9828 29374
rect 9884 28868 9940 29486
rect 10108 29428 10164 29438
rect 10332 29428 10388 30380
rect 10444 30322 10500 30334
rect 10444 30270 10446 30322
rect 10498 30270 10500 30322
rect 10444 30212 10500 30270
rect 10444 30146 10500 30156
rect 11004 30212 11060 30942
rect 11228 30660 11284 33852
rect 11340 33348 11396 33964
rect 11452 33954 11508 33964
rect 12012 34020 12068 34078
rect 12012 33954 12068 33964
rect 12124 33570 12180 33582
rect 12124 33518 12126 33570
rect 12178 33518 12180 33570
rect 11452 33348 11508 33358
rect 11340 33346 11508 33348
rect 11340 33294 11454 33346
rect 11506 33294 11508 33346
rect 11340 33292 11508 33294
rect 11452 33282 11508 33292
rect 11676 33346 11732 33358
rect 11676 33294 11678 33346
rect 11730 33294 11732 33346
rect 11676 33124 11732 33294
rect 11676 33058 11732 33068
rect 11452 32676 11508 32686
rect 11452 32452 11508 32620
rect 11452 32450 11732 32452
rect 11452 32398 11454 32450
rect 11506 32398 11732 32450
rect 11452 32396 11732 32398
rect 11452 32386 11508 32396
rect 11452 31666 11508 31678
rect 11452 31614 11454 31666
rect 11506 31614 11508 31666
rect 11228 30594 11284 30604
rect 11340 30994 11396 31006
rect 11340 30942 11342 30994
rect 11394 30942 11396 30994
rect 11004 30146 11060 30156
rect 10556 30100 10612 30110
rect 10556 30098 10948 30100
rect 10556 30046 10558 30098
rect 10610 30046 10948 30098
rect 10556 30044 10948 30046
rect 10556 30034 10612 30044
rect 10444 29652 10500 29662
rect 10444 29558 10500 29596
rect 10892 29650 10948 30044
rect 10892 29598 10894 29650
rect 10946 29598 10948 29650
rect 10892 29586 10948 29598
rect 10108 29334 10164 29372
rect 10220 29372 10388 29428
rect 10556 29428 10612 29438
rect 9884 28802 9940 28812
rect 10220 28980 10276 29372
rect 10556 29334 10612 29372
rect 9772 28690 9828 28700
rect 10108 28756 10164 28766
rect 10108 28662 10164 28700
rect 9660 28530 9716 28542
rect 9660 28478 9662 28530
rect 9714 28478 9716 28530
rect 9660 28084 9716 28478
rect 9660 28018 9716 28028
rect 10220 27858 10276 28924
rect 11004 29314 11060 29326
rect 11004 29262 11006 29314
rect 11058 29262 11060 29314
rect 10556 28868 10612 28878
rect 10444 28812 10556 28868
rect 10444 28642 10500 28812
rect 10556 28802 10612 28812
rect 11004 28756 11060 29262
rect 11340 28868 11396 30942
rect 11452 30996 11508 31614
rect 11564 31668 11620 31678
rect 11564 31574 11620 31612
rect 11452 30324 11508 30940
rect 11452 30258 11508 30268
rect 11340 28802 11396 28812
rect 11004 28690 11060 28700
rect 10444 28590 10446 28642
rect 10498 28590 10500 28642
rect 10444 28578 10500 28590
rect 10556 28644 10612 28654
rect 10444 28196 10500 28206
rect 10332 28084 10388 28094
rect 10332 27990 10388 28028
rect 10444 28082 10500 28140
rect 10444 28030 10446 28082
rect 10498 28030 10500 28082
rect 10444 28018 10500 28030
rect 10556 28082 10612 28588
rect 11452 28644 11508 28654
rect 11452 28550 11508 28588
rect 11004 28532 11060 28542
rect 10892 28530 11060 28532
rect 10892 28478 11006 28530
rect 11058 28478 11060 28530
rect 10892 28476 11060 28478
rect 10780 28420 10836 28430
rect 10556 28030 10558 28082
rect 10610 28030 10612 28082
rect 10556 28018 10612 28030
rect 10668 28364 10780 28420
rect 10220 27806 10222 27858
rect 10274 27806 10276 27858
rect 10220 27794 10276 27806
rect 9212 27234 9268 27244
rect 9884 27300 9940 27310
rect 8428 26962 8484 26984
rect 8428 26910 8430 26962
rect 8482 26910 8484 26962
rect 8428 26908 8484 26910
rect 8540 26908 8596 27132
rect 8316 26852 8596 26908
rect 7308 26572 7812 26628
rect 7308 25618 7364 26572
rect 7756 26514 7812 26572
rect 7756 26462 7758 26514
rect 7810 26462 7812 26514
rect 7756 26450 7812 26462
rect 7308 25566 7310 25618
rect 7362 25566 7364 25618
rect 7308 25554 7364 25566
rect 7532 26404 7588 26414
rect 6860 24946 7140 24948
rect 6860 24894 6862 24946
rect 6914 24894 7140 24946
rect 6860 24892 7140 24894
rect 6860 24724 6916 24892
rect 6860 24658 6916 24668
rect 7084 24052 7140 24062
rect 7084 23938 7140 23996
rect 7084 23886 7086 23938
rect 7138 23886 7140 23938
rect 7084 23874 7140 23886
rect 7196 23940 7252 23950
rect 7196 23846 7252 23884
rect 7308 23266 7364 23278
rect 7308 23214 7310 23266
rect 7362 23214 7364 23266
rect 7308 23156 7364 23214
rect 7364 23100 7476 23156
rect 7308 23090 7364 23100
rect 7196 22484 7252 22494
rect 6748 22430 6750 22482
rect 6802 22430 6804 22482
rect 6412 22372 6468 22382
rect 6188 22258 6244 22270
rect 6188 22206 6190 22258
rect 6242 22206 6244 22258
rect 6188 22148 6244 22206
rect 6188 22082 6244 22092
rect 6300 22146 6356 22158
rect 6300 22094 6302 22146
rect 6354 22094 6356 22146
rect 6188 21700 6244 21710
rect 6188 21586 6244 21644
rect 6188 21534 6190 21586
rect 6242 21534 6244 21586
rect 6188 21522 6244 21534
rect 6300 21140 6356 22094
rect 5964 20738 6020 20748
rect 6076 21084 6356 21140
rect 5516 20524 5796 20580
rect 5964 20578 6020 20590
rect 5964 20526 5966 20578
rect 6018 20526 6020 20578
rect 5180 20132 5236 20142
rect 5180 20038 5236 20076
rect 5516 19572 5572 20524
rect 5964 20468 6020 20526
rect 6076 20580 6132 21084
rect 6300 20916 6356 20926
rect 6412 20916 6468 22316
rect 6524 22148 6580 22158
rect 6524 21586 6580 22092
rect 6748 21812 6804 22430
rect 6748 21746 6804 21756
rect 7084 22482 7252 22484
rect 7084 22430 7198 22482
rect 7250 22430 7252 22482
rect 7084 22428 7252 22430
rect 6524 21534 6526 21586
rect 6578 21534 6580 21586
rect 6524 21522 6580 21534
rect 6636 21700 6692 21710
rect 6300 20914 6468 20916
rect 6300 20862 6302 20914
rect 6354 20862 6468 20914
rect 6300 20860 6468 20862
rect 6300 20850 6356 20860
rect 6188 20804 6244 20814
rect 6188 20710 6244 20748
rect 6524 20804 6580 20814
rect 6076 20524 6244 20580
rect 5628 20412 6020 20468
rect 5628 20132 5684 20412
rect 6076 20356 6132 20366
rect 5740 20300 6076 20356
rect 5740 20242 5796 20300
rect 6076 20290 6132 20300
rect 5740 20190 5742 20242
rect 5794 20190 5796 20242
rect 5740 20178 5796 20190
rect 5628 20038 5684 20076
rect 6188 20018 6244 20524
rect 6412 20578 6468 20590
rect 6412 20526 6414 20578
rect 6466 20526 6468 20578
rect 6412 20356 6468 20526
rect 6412 20290 6468 20300
rect 6412 20132 6468 20142
rect 6524 20132 6580 20748
rect 6412 20130 6580 20132
rect 6412 20078 6414 20130
rect 6466 20078 6580 20130
rect 6412 20076 6580 20078
rect 6636 20692 6692 21644
rect 6412 20066 6468 20076
rect 6188 19966 6190 20018
rect 6242 19966 6244 20018
rect 6188 19954 6244 19966
rect 6524 19908 6580 19918
rect 6636 19908 6692 20636
rect 6524 19906 6692 19908
rect 6524 19854 6526 19906
rect 6578 19854 6692 19906
rect 6524 19852 6692 19854
rect 6748 20802 6804 20814
rect 6748 20750 6750 20802
rect 6802 20750 6804 20802
rect 6524 19842 6580 19852
rect 5852 19796 5908 19806
rect 5852 19794 6132 19796
rect 5852 19742 5854 19794
rect 5906 19742 6132 19794
rect 5852 19740 6132 19742
rect 5852 19730 5908 19740
rect 5516 19516 5908 19572
rect 5180 19236 5236 19246
rect 5516 19236 5572 19246
rect 5180 19234 5572 19236
rect 5180 19182 5182 19234
rect 5234 19182 5518 19234
rect 5570 19182 5572 19234
rect 5180 19180 5572 19182
rect 5180 19170 5236 19180
rect 5516 19170 5572 19180
rect 5740 19236 5796 19246
rect 5740 19122 5796 19180
rect 5852 19236 5908 19516
rect 5852 19234 6020 19236
rect 5852 19182 5854 19234
rect 5906 19182 6020 19234
rect 5852 19180 6020 19182
rect 5852 19170 5908 19180
rect 5740 19070 5742 19122
rect 5794 19070 5796 19122
rect 5628 18676 5684 18686
rect 5740 18676 5796 19070
rect 5628 18674 5796 18676
rect 5628 18622 5630 18674
rect 5682 18622 5796 18674
rect 5628 18620 5796 18622
rect 5628 18610 5684 18620
rect 5068 17726 5070 17778
rect 5122 17726 5124 17778
rect 4732 17668 4788 17678
rect 5068 17668 5124 17726
rect 5964 17780 6020 19180
rect 6076 18676 6132 19740
rect 6300 19236 6356 19246
rect 6188 18676 6244 18686
rect 6076 18620 6188 18676
rect 6188 18582 6244 18620
rect 6300 18562 6356 19180
rect 6300 18510 6302 18562
rect 6354 18510 6356 18562
rect 6300 18498 6356 18510
rect 6524 18452 6580 18462
rect 6188 17780 6244 17790
rect 5964 17778 6244 17780
rect 5964 17726 6190 17778
rect 6242 17726 6244 17778
rect 5964 17724 6244 17726
rect 6188 17714 6244 17724
rect 6524 17780 6580 18396
rect 6748 18228 6804 20750
rect 6972 20802 7028 20814
rect 6972 20750 6974 20802
rect 7026 20750 7028 20802
rect 6972 20132 7028 20750
rect 6860 19236 6916 19246
rect 6972 19236 7028 20076
rect 7084 19906 7140 22428
rect 7196 22418 7252 22428
rect 7308 22148 7364 22158
rect 7196 22146 7364 22148
rect 7196 22094 7310 22146
rect 7362 22094 7364 22146
rect 7196 22092 7364 22094
rect 7196 20804 7252 22092
rect 7308 22082 7364 22092
rect 7420 21364 7476 23100
rect 7532 22708 7588 26348
rect 8316 26404 8372 26852
rect 8316 26338 8372 26348
rect 8652 26402 8708 26414
rect 8652 26350 8654 26402
rect 8706 26350 8708 26402
rect 7980 26292 8036 26302
rect 7868 26180 7924 26190
rect 7868 26086 7924 26124
rect 7980 25956 8036 26236
rect 7868 25900 8036 25956
rect 8092 26290 8148 26302
rect 8540 26292 8596 26302
rect 8092 26238 8094 26290
rect 8146 26238 8148 26290
rect 7644 25284 7700 25294
rect 7644 24050 7700 25228
rect 7868 24612 7924 25900
rect 7980 25506 8036 25518
rect 7980 25454 7982 25506
rect 8034 25454 8036 25506
rect 7980 25172 8036 25454
rect 7980 25106 8036 25116
rect 7980 24836 8036 24846
rect 8092 24836 8148 26238
rect 8428 26290 8596 26292
rect 8428 26238 8542 26290
rect 8594 26238 8596 26290
rect 8428 26236 8596 26238
rect 8204 25508 8260 25518
rect 8428 25508 8484 26236
rect 8540 26226 8596 26236
rect 8652 25620 8708 26350
rect 9548 26404 9604 26414
rect 8876 26292 8932 26302
rect 8876 26290 9492 26292
rect 8876 26238 8878 26290
rect 8930 26238 9492 26290
rect 8876 26236 9492 26238
rect 8876 26226 8932 26236
rect 8764 25732 8820 25742
rect 8764 25638 8820 25676
rect 8204 25506 8484 25508
rect 8204 25454 8206 25506
rect 8258 25454 8484 25506
rect 8204 25452 8484 25454
rect 8540 25564 8708 25620
rect 8204 25442 8260 25452
rect 7980 24834 8148 24836
rect 7980 24782 7982 24834
rect 8034 24782 8148 24834
rect 7980 24780 8148 24782
rect 7980 24770 8036 24780
rect 7868 24556 8260 24612
rect 7644 23998 7646 24050
rect 7698 23998 7700 24050
rect 7644 23986 7700 23998
rect 8092 23938 8148 23950
rect 8092 23886 8094 23938
rect 8146 23886 8148 23938
rect 8092 23716 8148 23886
rect 8092 23650 8148 23660
rect 8092 23268 8148 23278
rect 7532 22652 7700 22708
rect 7532 22484 7588 22494
rect 7532 22390 7588 22428
rect 7196 20738 7252 20748
rect 7308 21308 7476 21364
rect 7308 20020 7364 21308
rect 7644 20804 7700 22652
rect 7980 22484 8036 22494
rect 7980 22390 8036 22428
rect 8092 22260 8148 23212
rect 7756 22258 8148 22260
rect 7756 22206 8094 22258
rect 8146 22206 8148 22258
rect 7756 22204 8148 22206
rect 7756 21698 7812 22204
rect 8092 22036 8148 22204
rect 8204 22036 8260 24556
rect 8316 24500 8372 25452
rect 8540 25172 8596 25564
rect 9436 25506 9492 26236
rect 9436 25454 9438 25506
rect 9490 25454 9492 25506
rect 9436 25442 9492 25454
rect 9548 25732 9604 26348
rect 9660 26292 9716 26302
rect 9660 26198 9716 26236
rect 8652 25394 8708 25406
rect 8652 25342 8654 25394
rect 8706 25342 8708 25394
rect 8652 25284 8708 25342
rect 9548 25394 9604 25676
rect 9772 25508 9828 25518
rect 9772 25414 9828 25452
rect 9548 25342 9550 25394
rect 9602 25342 9604 25394
rect 9548 25330 9604 25342
rect 8652 25218 8708 25228
rect 8764 25282 8820 25294
rect 8764 25230 8766 25282
rect 8818 25230 8820 25282
rect 8428 25060 8484 25070
rect 8428 24722 8484 25004
rect 8428 24670 8430 24722
rect 8482 24670 8484 24722
rect 8428 24658 8484 24670
rect 8316 24444 8484 24500
rect 8316 23268 8372 23278
rect 8428 23268 8484 24444
rect 8540 24052 8596 25116
rect 8540 23958 8596 23996
rect 8764 23716 8820 25230
rect 9548 25060 9604 25070
rect 9548 24836 9604 25004
rect 9212 24834 9604 24836
rect 9212 24782 9550 24834
rect 9602 24782 9604 24834
rect 9212 24780 9604 24782
rect 8988 24724 9044 24734
rect 8876 24612 8932 24622
rect 8988 24612 9044 24668
rect 8876 24610 9044 24612
rect 8876 24558 8878 24610
rect 8930 24558 9044 24610
rect 8876 24556 9044 24558
rect 8876 24546 8932 24556
rect 8764 23650 8820 23660
rect 8652 23268 8708 23278
rect 8428 23266 8708 23268
rect 8428 23214 8654 23266
rect 8706 23214 8708 23266
rect 8428 23212 8708 23214
rect 8316 23154 8372 23212
rect 8652 23202 8708 23212
rect 8316 23102 8318 23154
rect 8370 23102 8372 23154
rect 8316 23090 8372 23102
rect 8764 23154 8820 23166
rect 8764 23102 8766 23154
rect 8818 23102 8820 23154
rect 8428 23042 8484 23054
rect 8428 22990 8430 23042
rect 8482 22990 8484 23042
rect 8428 22596 8484 22990
rect 8652 22820 8708 22830
rect 8316 22370 8372 22382
rect 8316 22318 8318 22370
rect 8370 22318 8372 22370
rect 8316 22260 8372 22318
rect 8428 22260 8484 22540
rect 8316 22204 8428 22260
rect 8428 22194 8484 22204
rect 8540 22764 8652 22820
rect 8204 21980 8372 22036
rect 8092 21970 8148 21980
rect 7756 21646 7758 21698
rect 7810 21646 7812 21698
rect 7756 21634 7812 21646
rect 8092 21588 8148 21598
rect 7980 21586 8148 21588
rect 7980 21534 8094 21586
rect 8146 21534 8148 21586
rect 7980 21532 8148 21534
rect 7980 20914 8036 21532
rect 8092 21522 8148 21532
rect 8316 21586 8372 21980
rect 8540 21810 8596 22764
rect 8652 22754 8708 22764
rect 8652 22484 8708 22494
rect 8652 22390 8708 22428
rect 8764 22372 8820 23102
rect 8764 22306 8820 22316
rect 8540 21758 8542 21810
rect 8594 21758 8596 21810
rect 8540 21746 8596 21758
rect 8764 22146 8820 22158
rect 8764 22094 8766 22146
rect 8818 22094 8820 22146
rect 8764 21698 8820 22094
rect 8876 22148 8932 22158
rect 8988 22148 9044 24556
rect 9212 24162 9268 24780
rect 9548 24770 9604 24780
rect 9660 24500 9716 24510
rect 9660 24498 9828 24500
rect 9660 24446 9662 24498
rect 9714 24446 9828 24498
rect 9660 24444 9828 24446
rect 9660 24434 9716 24444
rect 9212 24110 9214 24162
rect 9266 24110 9268 24162
rect 9212 24098 9268 24110
rect 9548 24050 9604 24062
rect 9548 23998 9550 24050
rect 9602 23998 9604 24050
rect 9436 23828 9492 23838
rect 9436 23734 9492 23772
rect 9548 23492 9604 23998
rect 9548 23426 9604 23436
rect 9772 23716 9828 24444
rect 9660 23268 9716 23278
rect 9660 23174 9716 23212
rect 9548 23156 9604 23166
rect 9548 23062 9604 23100
rect 9772 22932 9828 23660
rect 9772 22866 9828 22876
rect 9212 22820 9268 22830
rect 9212 22370 9268 22764
rect 9884 22708 9940 27244
rect 10444 27300 10500 27310
rect 10444 27206 10500 27244
rect 10668 26962 10724 28364
rect 10780 28354 10836 28364
rect 10780 27860 10836 27870
rect 10892 27860 10948 28476
rect 11004 28466 11060 28476
rect 10780 27858 10948 27860
rect 10780 27806 10782 27858
rect 10834 27806 10948 27858
rect 10780 27804 10948 27806
rect 10780 27794 10836 27804
rect 11452 27746 11508 27758
rect 11452 27694 11454 27746
rect 11506 27694 11508 27746
rect 10668 26910 10670 26962
rect 10722 26910 10724 26962
rect 10668 26908 10724 26910
rect 10220 26852 10724 26908
rect 10780 27186 10836 27198
rect 10780 27134 10782 27186
rect 10834 27134 10836 27186
rect 10780 26908 10836 27134
rect 11116 26962 11172 26974
rect 11116 26910 11118 26962
rect 11170 26910 11172 26962
rect 10780 26852 11060 26908
rect 10220 26850 10276 26852
rect 10220 26798 10222 26850
rect 10274 26798 10276 26850
rect 10220 26786 10276 26798
rect 11004 26180 11060 26852
rect 11116 26404 11172 26910
rect 11228 26962 11284 26974
rect 11228 26910 11230 26962
rect 11282 26910 11284 26962
rect 11228 26516 11284 26910
rect 11452 26964 11508 27694
rect 11452 26898 11508 26908
rect 11228 26450 11284 26460
rect 11340 26850 11396 26862
rect 11340 26798 11342 26850
rect 11394 26798 11396 26850
rect 11116 26338 11172 26348
rect 11340 26404 11396 26798
rect 11340 26338 11396 26348
rect 11004 26124 11620 26180
rect 10444 25618 10500 25630
rect 10444 25566 10446 25618
rect 10498 25566 10500 25618
rect 10332 25506 10388 25518
rect 10332 25454 10334 25506
rect 10386 25454 10388 25506
rect 10108 25060 10164 25070
rect 10108 24946 10164 25004
rect 10108 24894 10110 24946
rect 10162 24894 10164 24946
rect 10108 24882 10164 24894
rect 10220 24948 10276 24958
rect 10220 24854 10276 24892
rect 9996 24724 10052 24762
rect 9996 24658 10052 24668
rect 9660 22652 9940 22708
rect 9996 24500 10052 24510
rect 9324 22596 9380 22606
rect 9324 22484 9380 22540
rect 9324 22428 9492 22484
rect 9212 22318 9214 22370
rect 9266 22318 9268 22370
rect 9212 22306 9268 22318
rect 9436 22372 9492 22428
rect 9436 22316 9604 22372
rect 9548 22258 9604 22316
rect 9548 22206 9550 22258
rect 9602 22206 9604 22258
rect 9548 22194 9604 22206
rect 8988 22092 9380 22148
rect 8876 22054 8932 22092
rect 8764 21646 8766 21698
rect 8818 21646 8820 21698
rect 8764 21634 8820 21646
rect 8316 21534 8318 21586
rect 8370 21534 8372 21586
rect 8204 21474 8260 21486
rect 8204 21422 8206 21474
rect 8258 21422 8260 21474
rect 8204 21028 8260 21422
rect 8316 21140 8372 21534
rect 8316 21084 8596 21140
rect 8204 20962 8260 20972
rect 7980 20862 7982 20914
rect 8034 20862 8036 20914
rect 7980 20850 8036 20862
rect 7644 20748 7924 20804
rect 7420 20692 7476 20702
rect 7868 20692 7924 20748
rect 8428 20802 8484 20814
rect 8428 20750 8430 20802
rect 8482 20750 8484 20802
rect 8428 20692 8484 20750
rect 7868 20636 8260 20692
rect 7420 20598 7476 20636
rect 7532 20578 7588 20590
rect 7532 20526 7534 20578
rect 7586 20526 7588 20578
rect 7308 20018 7476 20020
rect 7308 19966 7310 20018
rect 7362 19966 7476 20018
rect 7308 19964 7476 19966
rect 7308 19954 7364 19964
rect 7084 19854 7086 19906
rect 7138 19854 7140 19906
rect 7084 19842 7140 19854
rect 6860 19234 7028 19236
rect 6860 19182 6862 19234
rect 6914 19182 7028 19234
rect 6860 19180 7028 19182
rect 7420 19236 7476 19964
rect 7532 19460 7588 20526
rect 7644 20578 7700 20590
rect 7644 20526 7646 20578
rect 7698 20526 7700 20578
rect 7644 20356 7700 20526
rect 7644 20290 7700 20300
rect 7644 20020 7700 20030
rect 7644 19684 7700 19964
rect 7868 20020 7924 20030
rect 7868 19926 7924 19964
rect 7644 19618 7700 19628
rect 7980 19908 8036 20636
rect 8204 20130 8260 20636
rect 8428 20626 8484 20636
rect 8204 20078 8206 20130
rect 8258 20078 8260 20130
rect 8204 20066 8260 20078
rect 8316 20132 8372 20142
rect 7532 19394 7588 19404
rect 7756 19346 7812 19358
rect 7756 19294 7758 19346
rect 7810 19294 7812 19346
rect 7756 19236 7812 19294
rect 7420 19180 7812 19236
rect 6860 19170 6916 19180
rect 6860 18676 6916 18686
rect 6860 18562 6916 18620
rect 6860 18510 6862 18562
rect 6914 18510 6916 18562
rect 6860 18498 6916 18510
rect 6972 18564 7028 19180
rect 7980 18676 8036 19852
rect 8316 19346 8372 20076
rect 8428 20020 8484 20030
rect 8540 20020 8596 21084
rect 8876 20802 8932 20814
rect 8876 20750 8878 20802
rect 8930 20750 8932 20802
rect 8876 20356 8932 20750
rect 8876 20290 8932 20300
rect 9212 20692 9268 20702
rect 9324 20692 9380 22092
rect 9436 22146 9492 22158
rect 9436 22094 9438 22146
rect 9490 22094 9492 22146
rect 9436 22036 9492 22094
rect 9436 21970 9492 21980
rect 9548 21812 9604 21822
rect 9660 21812 9716 22652
rect 9996 22594 10052 24444
rect 10332 23938 10388 25454
rect 10444 25508 10500 25566
rect 10444 25442 10500 25452
rect 11564 25506 11620 26124
rect 11564 25454 11566 25506
rect 11618 25454 11620 25506
rect 11564 25442 11620 25454
rect 11228 25396 11284 25406
rect 11228 25302 11284 25340
rect 10332 23886 10334 23938
rect 10386 23886 10388 23938
rect 10220 23492 10276 23502
rect 10220 23044 10276 23436
rect 10332 23268 10388 23886
rect 10444 24834 10500 24846
rect 10444 24782 10446 24834
rect 10498 24782 10500 24834
rect 10444 23828 10500 24782
rect 10668 24836 10724 24846
rect 10668 24050 10724 24780
rect 11340 24836 11396 24846
rect 11340 24742 11396 24780
rect 11228 24722 11284 24734
rect 11228 24670 11230 24722
rect 11282 24670 11284 24722
rect 11228 24500 11284 24670
rect 11228 24434 11284 24444
rect 10668 23998 10670 24050
rect 10722 23998 10724 24050
rect 10668 23986 10724 23998
rect 10556 23940 10612 23950
rect 10556 23846 10612 23884
rect 11564 23940 11620 23950
rect 10444 23762 10500 23772
rect 11116 23826 11172 23838
rect 11116 23774 11118 23826
rect 11170 23774 11172 23826
rect 10332 23202 10388 23212
rect 11116 23268 11172 23774
rect 11116 23202 11172 23212
rect 11564 23154 11620 23884
rect 11676 23492 11732 32396
rect 12124 31668 12180 33518
rect 12236 32900 12292 35308
rect 12348 35698 12404 35710
rect 12348 35646 12350 35698
rect 12402 35646 12404 35698
rect 12348 35028 12404 35646
rect 12460 35028 12516 35038
rect 12348 34972 12460 35028
rect 12460 34934 12516 34972
rect 12684 34132 12740 34142
rect 12684 34038 12740 34076
rect 12796 34020 12852 34030
rect 12236 32844 12628 32900
rect 12572 32788 12628 32844
rect 12572 32674 12628 32732
rect 12572 32622 12574 32674
rect 12626 32622 12628 32674
rect 12572 32610 12628 32622
rect 12796 32676 12852 33964
rect 12796 32562 12852 32620
rect 12796 32510 12798 32562
rect 12850 32510 12852 32562
rect 12796 32498 12852 32510
rect 12012 31612 12124 31668
rect 11788 31554 11844 31566
rect 11788 31502 11790 31554
rect 11842 31502 11844 31554
rect 11788 30772 11844 31502
rect 11788 30706 11844 30716
rect 11900 30212 11956 30222
rect 11900 30118 11956 30156
rect 12012 30098 12068 31612
rect 12124 31602 12180 31612
rect 12572 32116 12628 32126
rect 12124 30996 12180 31006
rect 12124 30902 12180 30940
rect 12460 30772 12516 30782
rect 12236 30212 12292 30222
rect 12236 30118 12292 30156
rect 12460 30210 12516 30716
rect 12460 30158 12462 30210
rect 12514 30158 12516 30210
rect 12460 30146 12516 30158
rect 12012 30046 12014 30098
rect 12066 30046 12068 30098
rect 12012 30034 12068 30046
rect 12572 30098 12628 32060
rect 12796 30884 12852 30894
rect 12796 30210 12852 30828
rect 12796 30158 12798 30210
rect 12850 30158 12852 30210
rect 12796 30146 12852 30158
rect 12572 30046 12574 30098
rect 12626 30046 12628 30098
rect 12572 30034 12628 30046
rect 11900 28980 11956 28990
rect 11788 28866 11844 28878
rect 11788 28814 11790 28866
rect 11842 28814 11844 28866
rect 11788 27858 11844 28814
rect 11900 28754 11956 28924
rect 11900 28702 11902 28754
rect 11954 28702 11956 28754
rect 11900 28690 11956 28702
rect 12908 28866 12964 35868
rect 13132 35858 13188 35868
rect 13580 35924 13636 36540
rect 13804 36372 13860 36382
rect 14588 36372 14644 36382
rect 13804 36370 14644 36372
rect 13804 36318 13806 36370
rect 13858 36318 14590 36370
rect 14642 36318 14644 36370
rect 13804 36316 14644 36318
rect 13804 36306 13860 36316
rect 14588 36306 14644 36316
rect 14700 36148 14756 37436
rect 14812 37044 14868 37774
rect 15260 37826 15316 37838
rect 15260 37774 15262 37826
rect 15314 37774 15316 37826
rect 14812 36978 14868 36988
rect 15148 37042 15204 37054
rect 15148 36990 15150 37042
rect 15202 36990 15204 37042
rect 15148 36932 15204 36990
rect 14924 36876 15148 36932
rect 14924 36706 14980 36876
rect 15148 36866 15204 36876
rect 14924 36654 14926 36706
rect 14978 36654 14980 36706
rect 14924 36642 14980 36654
rect 15260 36484 15316 37774
rect 15932 37828 15988 38558
rect 15932 37490 15988 37772
rect 15932 37438 15934 37490
rect 15986 37438 15988 37490
rect 15932 37426 15988 37438
rect 16156 37492 16212 41200
rect 16828 38668 16884 41200
rect 16716 38612 16884 38668
rect 16716 38610 16772 38612
rect 16716 38558 16718 38610
rect 16770 38558 16772 38610
rect 16716 38546 16772 38558
rect 16716 38388 16772 38398
rect 16156 37426 16212 37436
rect 16268 37826 16324 37838
rect 16268 37774 16270 37826
rect 16322 37774 16324 37826
rect 16268 37268 16324 37774
rect 16156 37212 16324 37268
rect 16716 37266 16772 38332
rect 17500 38388 17556 41200
rect 18172 38668 18228 41200
rect 18844 38668 18900 41200
rect 18172 38612 18340 38668
rect 17500 38322 17556 38332
rect 18172 38276 18228 38286
rect 18172 38182 18228 38220
rect 17500 38050 17556 38062
rect 17500 37998 17502 38050
rect 17554 37998 17556 38050
rect 16716 37214 16718 37266
rect 16770 37214 16772 37266
rect 15484 37156 15540 37166
rect 15484 37154 15652 37156
rect 15484 37102 15486 37154
rect 15538 37102 15652 37154
rect 15484 37100 15652 37102
rect 15484 37090 15540 37100
rect 15260 36418 15316 36428
rect 15372 37044 15428 37054
rect 15372 36482 15428 36988
rect 15372 36430 15374 36482
rect 15426 36430 15428 36482
rect 15372 36418 15428 36430
rect 14028 36092 14756 36148
rect 13916 36036 13972 36046
rect 13916 35924 13972 35980
rect 13580 35922 13972 35924
rect 13580 35870 13582 35922
rect 13634 35870 13972 35922
rect 13580 35868 13972 35870
rect 13580 35858 13636 35868
rect 13916 35810 13972 35868
rect 14028 35922 14084 36092
rect 14028 35870 14030 35922
rect 14082 35870 14084 35922
rect 14028 35858 14084 35870
rect 14588 35868 14868 35924
rect 13916 35758 13918 35810
rect 13970 35758 13972 35810
rect 13916 35746 13972 35758
rect 14476 35810 14532 35822
rect 14476 35758 14478 35810
rect 14530 35758 14532 35810
rect 14364 35698 14420 35710
rect 14364 35646 14366 35698
rect 14418 35646 14420 35698
rect 13916 35588 13972 35598
rect 13916 34804 13972 35532
rect 14364 35308 14420 35646
rect 14476 35588 14532 35758
rect 14476 35522 14532 35532
rect 14140 35252 14420 35308
rect 14028 34916 14084 34926
rect 14028 34822 14084 34860
rect 13804 34802 13972 34804
rect 13804 34750 13918 34802
rect 13970 34750 13972 34802
rect 13804 34748 13972 34750
rect 13020 34692 13076 34702
rect 13020 34598 13076 34636
rect 13692 34692 13748 34702
rect 13692 33572 13748 34636
rect 13692 33506 13748 33516
rect 13804 33348 13860 34748
rect 13916 34738 13972 34748
rect 14140 34802 14196 35252
rect 14476 34916 14532 34926
rect 14588 34916 14644 35868
rect 14812 35812 14868 35868
rect 14924 35812 14980 35822
rect 15148 35812 15204 35822
rect 14812 35810 14980 35812
rect 14812 35758 14926 35810
rect 14978 35758 14980 35810
rect 14812 35756 14980 35758
rect 14924 35746 14980 35756
rect 15036 35810 15204 35812
rect 15036 35758 15150 35810
rect 15202 35758 15204 35810
rect 15036 35756 15204 35758
rect 14532 34860 14644 34916
rect 14700 35698 14756 35710
rect 14700 35646 14702 35698
rect 14754 35646 14756 35698
rect 14700 34916 14756 35646
rect 15036 35476 15092 35756
rect 15148 35746 15204 35756
rect 15036 35410 15092 35420
rect 15148 35586 15204 35598
rect 15596 35588 15652 37100
rect 15708 37044 15764 37054
rect 15764 36988 15876 37044
rect 15708 36978 15764 36988
rect 15708 36370 15764 36382
rect 15708 36318 15710 36370
rect 15762 36318 15764 36370
rect 15708 36260 15764 36318
rect 15708 36194 15764 36204
rect 15708 35812 15764 35822
rect 15708 35718 15764 35756
rect 15148 35534 15150 35586
rect 15202 35534 15204 35586
rect 14924 35140 14980 35150
rect 14476 34822 14532 34860
rect 14700 34850 14756 34860
rect 14812 35026 14868 35038
rect 14812 34974 14814 35026
rect 14866 34974 14868 35026
rect 14140 34750 14142 34802
rect 14194 34750 14196 34802
rect 13916 34242 13972 34254
rect 13916 34190 13918 34242
rect 13970 34190 13972 34242
rect 13916 34132 13972 34190
rect 13916 34066 13972 34076
rect 14028 34130 14084 34142
rect 14028 34078 14030 34130
rect 14082 34078 14084 34130
rect 13804 33282 13860 33292
rect 13916 33906 13972 33918
rect 13916 33854 13918 33906
rect 13970 33854 13972 33906
rect 13692 33236 13748 33246
rect 13580 32788 13636 32798
rect 13580 32694 13636 32732
rect 13692 32676 13748 33180
rect 13692 32582 13748 32620
rect 13132 32340 13188 32350
rect 13132 32338 13412 32340
rect 13132 32286 13134 32338
rect 13186 32286 13412 32338
rect 13132 32284 13412 32286
rect 13132 32274 13188 32284
rect 13356 31892 13412 32284
rect 13580 32338 13636 32350
rect 13580 32286 13582 32338
rect 13634 32286 13636 32338
rect 13468 32116 13524 32126
rect 13580 32116 13636 32286
rect 13524 32060 13636 32116
rect 13468 32050 13524 32060
rect 13916 31892 13972 33854
rect 14028 33796 14084 34078
rect 14140 33908 14196 34750
rect 14812 34804 14868 34974
rect 14812 34738 14868 34748
rect 14700 34692 14756 34730
rect 14700 34626 14756 34636
rect 14476 34580 14532 34590
rect 14476 34354 14532 34524
rect 14476 34302 14478 34354
rect 14530 34302 14532 34354
rect 14476 34290 14532 34302
rect 14700 34468 14756 34478
rect 14700 34354 14756 34412
rect 14700 34302 14702 34354
rect 14754 34302 14756 34354
rect 14700 34290 14756 34302
rect 14924 34354 14980 35084
rect 14924 34302 14926 34354
rect 14978 34302 14980 34354
rect 14924 34290 14980 34302
rect 15036 34132 15092 34142
rect 15148 34132 15204 35534
rect 15372 35532 15652 35588
rect 15708 35586 15764 35598
rect 15708 35534 15710 35586
rect 15762 35534 15764 35586
rect 15260 35476 15316 35486
rect 15260 35140 15316 35420
rect 15372 35140 15428 35532
rect 15708 35476 15764 35534
rect 15708 35410 15764 35420
rect 15484 35140 15540 35150
rect 15372 35138 15764 35140
rect 15372 35086 15486 35138
rect 15538 35086 15764 35138
rect 15372 35084 15764 35086
rect 15260 35074 15316 35084
rect 15484 35074 15540 35084
rect 15260 34692 15316 34702
rect 15260 34468 15316 34636
rect 15372 34690 15428 34702
rect 15372 34638 15374 34690
rect 15426 34638 15428 34690
rect 15372 34580 15428 34638
rect 15372 34524 15652 34580
rect 15596 34468 15652 34524
rect 15260 34412 15540 34468
rect 15372 34132 15428 34142
rect 15148 34130 15428 34132
rect 15148 34078 15374 34130
rect 15426 34078 15428 34130
rect 15148 34076 15428 34078
rect 14812 34020 14868 34030
rect 14812 34018 14980 34020
rect 14812 33966 14814 34018
rect 14866 33966 14980 34018
rect 14812 33964 14980 33966
rect 14812 33954 14868 33964
rect 14140 33852 14420 33908
rect 14028 33730 14084 33740
rect 14140 32450 14196 32462
rect 14140 32398 14142 32450
rect 14194 32398 14196 32450
rect 13356 31836 13636 31892
rect 13580 31780 13636 31836
rect 13916 31826 13972 31836
rect 14028 32338 14084 32350
rect 14028 32286 14030 32338
rect 14082 32286 14084 32338
rect 13580 31778 13860 31780
rect 13580 31726 13582 31778
rect 13634 31726 13860 31778
rect 13580 31724 13860 31726
rect 13580 31714 13636 31724
rect 13020 31668 13076 31678
rect 13020 30994 13076 31612
rect 13468 31668 13524 31678
rect 13468 31574 13524 31612
rect 13692 31220 13748 31230
rect 13468 31108 13524 31118
rect 13468 31014 13524 31052
rect 13020 30942 13022 30994
rect 13074 30942 13076 30994
rect 13020 30930 13076 30942
rect 13692 30212 13748 31164
rect 13804 31106 13860 31724
rect 13804 31054 13806 31106
rect 13858 31054 13860 31106
rect 13804 31042 13860 31054
rect 13916 31668 13972 31678
rect 13916 30994 13972 31612
rect 14028 31108 14084 32286
rect 14140 32116 14196 32398
rect 14140 32050 14196 32060
rect 14364 31668 14420 33852
rect 14588 33796 14644 33806
rect 14588 33570 14644 33740
rect 14588 33518 14590 33570
rect 14642 33518 14644 33570
rect 14588 33506 14644 33518
rect 14700 33348 14756 33358
rect 14700 33254 14756 33292
rect 14924 32900 14980 33964
rect 15036 33458 15092 34076
rect 15372 34066 15428 34076
rect 15036 33406 15038 33458
rect 15090 33406 15092 33458
rect 15036 33394 15092 33406
rect 15484 33346 15540 34412
rect 15596 34402 15652 34412
rect 15708 34244 15764 35084
rect 15820 35028 15876 36988
rect 16156 36932 16212 37212
rect 16716 37202 16772 37214
rect 17164 37826 17220 37838
rect 17164 37774 17166 37826
rect 17218 37774 17220 37826
rect 16156 36594 16212 36876
rect 16156 36542 16158 36594
rect 16210 36542 16212 36594
rect 16156 36530 16212 36542
rect 16380 37154 16436 37166
rect 16380 37102 16382 37154
rect 16434 37102 16436 37154
rect 16268 36258 16324 36270
rect 16268 36206 16270 36258
rect 16322 36206 16324 36258
rect 15932 36148 15988 36158
rect 16268 36148 16324 36206
rect 15932 35810 15988 36092
rect 15932 35758 15934 35810
rect 15986 35758 15988 35810
rect 15932 35746 15988 35758
rect 16044 36092 16324 36148
rect 16380 36148 16436 37102
rect 16492 36484 16548 36494
rect 17052 36484 17108 36494
rect 16492 36390 16548 36428
rect 16604 36482 17108 36484
rect 16604 36430 17054 36482
rect 17106 36430 17108 36482
rect 16604 36428 17108 36430
rect 16044 35252 16100 36092
rect 16380 36082 16436 36092
rect 16604 36036 16660 36428
rect 17052 36418 17108 36428
rect 16492 35980 16660 36036
rect 16716 36260 16772 36270
rect 16492 35924 16548 35980
rect 16380 35868 16548 35924
rect 16380 35810 16436 35868
rect 16380 35758 16382 35810
rect 16434 35758 16436 35810
rect 16380 35746 16436 35758
rect 16044 35186 16100 35196
rect 16268 35698 16324 35710
rect 16268 35646 16270 35698
rect 16322 35646 16324 35698
rect 15820 34972 15988 35028
rect 15820 34804 15876 34814
rect 15820 34710 15876 34748
rect 15596 34132 15652 34142
rect 15596 34038 15652 34076
rect 15708 33460 15764 34188
rect 15820 33460 15876 33470
rect 15708 33458 15876 33460
rect 15708 33406 15822 33458
rect 15874 33406 15876 33458
rect 15708 33404 15876 33406
rect 15820 33394 15876 33404
rect 15484 33294 15486 33346
rect 15538 33294 15540 33346
rect 15484 33282 15540 33294
rect 14924 32844 15204 32900
rect 14700 32562 14756 32574
rect 14700 32510 14702 32562
rect 14754 32510 14756 32562
rect 14700 32004 14756 32510
rect 14924 32562 14980 32574
rect 14924 32510 14926 32562
rect 14978 32510 14980 32562
rect 14364 31602 14420 31612
rect 14476 31948 14756 32004
rect 14812 32450 14868 32462
rect 14812 32398 14814 32450
rect 14866 32398 14868 32450
rect 14028 31042 14084 31052
rect 13916 30942 13918 30994
rect 13970 30942 13972 30994
rect 13916 30930 13972 30942
rect 14252 30884 14308 30894
rect 14476 30884 14532 31948
rect 14700 31780 14756 31790
rect 14700 31218 14756 31724
rect 14700 31166 14702 31218
rect 14754 31166 14756 31218
rect 14700 31154 14756 31166
rect 14812 31108 14868 32398
rect 14924 31892 14980 32510
rect 14924 31220 14980 31836
rect 14924 31154 14980 31164
rect 14812 31042 14868 31052
rect 15036 30994 15092 32844
rect 15148 32786 15204 32844
rect 15148 32734 15150 32786
rect 15202 32734 15204 32786
rect 15148 32722 15204 32734
rect 15036 30942 15038 30994
rect 15090 30942 15092 30994
rect 15036 30930 15092 30942
rect 15260 31778 15316 31790
rect 15260 31726 15262 31778
rect 15314 31726 15316 31778
rect 14252 30882 14532 30884
rect 14252 30830 14254 30882
rect 14306 30830 14532 30882
rect 14252 30828 14532 30830
rect 14588 30882 14644 30894
rect 14588 30830 14590 30882
rect 14642 30830 14644 30882
rect 14252 30818 14308 30828
rect 14588 30660 14644 30830
rect 15260 30884 15316 31726
rect 15596 31668 15652 31678
rect 15372 31220 15428 31230
rect 15372 31126 15428 31164
rect 15596 31218 15652 31612
rect 15596 31166 15598 31218
rect 15650 31166 15652 31218
rect 15596 31154 15652 31166
rect 15484 30996 15540 31006
rect 15260 30818 15316 30828
rect 15372 30940 15484 30996
rect 14140 30604 14644 30660
rect 14028 30324 14084 30334
rect 14140 30324 14196 30604
rect 14252 30436 14308 30446
rect 14252 30342 14308 30380
rect 14028 30322 14196 30324
rect 14028 30270 14030 30322
rect 14082 30270 14196 30322
rect 14028 30268 14196 30270
rect 15372 30322 15428 30940
rect 15484 30902 15540 30940
rect 15372 30270 15374 30322
rect 15426 30270 15428 30322
rect 13804 30212 13860 30222
rect 13692 30210 13860 30212
rect 13692 30158 13806 30210
rect 13858 30158 13860 30210
rect 13692 30156 13860 30158
rect 13804 30146 13860 30156
rect 14028 30212 14084 30268
rect 15372 30258 15428 30270
rect 14028 30146 14084 30156
rect 14476 30212 14532 30222
rect 14476 30118 14532 30156
rect 15484 30212 15540 30222
rect 14588 29988 14644 29998
rect 14924 29988 14980 29998
rect 14140 29876 14196 29886
rect 13692 29538 13748 29550
rect 13692 29486 13694 29538
rect 13746 29486 13748 29538
rect 12908 28814 12910 28866
rect 12962 28814 12964 28866
rect 12908 28754 12964 28814
rect 12908 28702 12910 28754
rect 12962 28702 12964 28754
rect 12460 28644 12516 28654
rect 11788 27806 11790 27858
rect 11842 27806 11844 27858
rect 11788 27794 11844 27806
rect 12236 27858 12292 27870
rect 12236 27806 12238 27858
rect 12290 27806 12292 27858
rect 12236 27186 12292 27806
rect 12236 27134 12238 27186
rect 12290 27134 12292 27186
rect 12236 27122 12292 27134
rect 12348 26964 12404 27002
rect 12348 26898 12404 26908
rect 12124 26850 12180 26862
rect 12124 26798 12126 26850
rect 12178 26798 12180 26850
rect 12124 25618 12180 26798
rect 12124 25566 12126 25618
rect 12178 25566 12180 25618
rect 12124 25554 12180 25566
rect 12012 25508 12068 25518
rect 12012 25414 12068 25452
rect 12460 25508 12516 28588
rect 12908 27748 12964 28702
rect 13580 29426 13636 29438
rect 13580 29374 13582 29426
rect 13634 29374 13636 29426
rect 13580 28642 13636 29374
rect 13580 28590 13582 28642
rect 13634 28590 13636 28642
rect 13580 28084 13636 28590
rect 13692 28530 13748 29486
rect 14140 28868 14196 29820
rect 14588 29650 14644 29932
rect 14588 29598 14590 29650
rect 14642 29598 14644 29650
rect 14588 29586 14644 29598
rect 14700 29986 14980 29988
rect 14700 29934 14926 29986
rect 14978 29934 14980 29986
rect 14700 29932 14980 29934
rect 14700 29426 14756 29932
rect 14924 29922 14980 29932
rect 15484 29538 15540 30156
rect 15484 29486 15486 29538
rect 15538 29486 15540 29538
rect 15484 29474 15540 29486
rect 14700 29374 14702 29426
rect 14754 29374 14756 29426
rect 14700 29362 14756 29374
rect 14140 28754 14196 28812
rect 14140 28702 14142 28754
rect 14194 28702 14196 28754
rect 14140 28690 14196 28702
rect 15484 28756 15540 28766
rect 15484 28662 15540 28700
rect 13692 28478 13694 28530
rect 13746 28478 13748 28530
rect 13692 28196 13748 28478
rect 14364 28644 14420 28654
rect 13692 28140 14196 28196
rect 13580 28028 13860 28084
rect 12908 27682 12964 27692
rect 13356 27748 13412 27758
rect 13356 27074 13412 27692
rect 13356 27022 13358 27074
rect 13410 27022 13412 27074
rect 12572 26852 12628 26862
rect 12572 26758 12628 26796
rect 12908 26516 12964 26526
rect 12684 26404 12740 26414
rect 12460 25442 12516 25452
rect 12572 25620 12628 25630
rect 12124 25396 12180 25406
rect 12124 25302 12180 25340
rect 11788 25282 11844 25294
rect 11788 25230 11790 25282
rect 11842 25230 11844 25282
rect 11788 25060 11844 25230
rect 11788 24994 11844 25004
rect 12012 23938 12068 23950
rect 12012 23886 12014 23938
rect 12066 23886 12068 23938
rect 12012 23828 12068 23886
rect 12572 23938 12628 25564
rect 12684 25618 12740 26348
rect 12684 25566 12686 25618
rect 12738 25566 12740 25618
rect 12684 25554 12740 25566
rect 12796 25284 12852 25294
rect 12796 25190 12852 25228
rect 12908 24722 12964 26460
rect 13356 26404 13412 27022
rect 13468 26852 13524 26862
rect 13524 26796 13636 26852
rect 13468 26786 13524 26796
rect 12908 24670 12910 24722
rect 12962 24670 12964 24722
rect 12908 24658 12964 24670
rect 13244 26402 13412 26404
rect 13244 26350 13358 26402
rect 13410 26350 13412 26402
rect 13244 26348 13412 26350
rect 13244 24052 13300 26348
rect 13356 26338 13412 26348
rect 13580 25730 13636 26796
rect 13580 25678 13582 25730
rect 13634 25678 13636 25730
rect 13580 25666 13636 25678
rect 13692 25732 13748 25742
rect 13356 25620 13412 25630
rect 13412 25564 13524 25620
rect 13356 25554 13412 25564
rect 13468 25508 13524 25564
rect 13468 25452 13636 25508
rect 13580 25394 13636 25452
rect 13692 25506 13748 25676
rect 13692 25454 13694 25506
rect 13746 25454 13748 25506
rect 13692 25442 13748 25454
rect 13580 25342 13582 25394
rect 13634 25342 13636 25394
rect 13580 25330 13636 25342
rect 13468 25284 13524 25294
rect 13468 24276 13524 25228
rect 13804 24946 13860 28028
rect 14028 27074 14084 27086
rect 14028 27022 14030 27074
rect 14082 27022 14084 27074
rect 14028 25394 14084 27022
rect 14028 25342 14030 25394
rect 14082 25342 14084 25394
rect 14028 25330 14084 25342
rect 13804 24894 13806 24946
rect 13858 24894 13860 24946
rect 13804 24882 13860 24894
rect 13468 24220 13748 24276
rect 13244 23986 13300 23996
rect 13692 24050 13748 24220
rect 13692 23998 13694 24050
rect 13746 23998 13748 24050
rect 12572 23886 12574 23938
rect 12626 23886 12628 23938
rect 12572 23874 12628 23886
rect 12012 23762 12068 23772
rect 13468 23828 13524 23838
rect 13468 23734 13524 23772
rect 13692 23716 13748 23998
rect 13692 23650 13748 23660
rect 11676 23426 11732 23436
rect 12124 23268 12180 23278
rect 12124 23174 12180 23212
rect 11564 23102 11566 23154
rect 11618 23102 11620 23154
rect 11564 23090 11620 23102
rect 10220 22988 10388 23044
rect 9996 22542 9998 22594
rect 10050 22542 10052 22594
rect 9996 22530 10052 22542
rect 10220 22372 10276 22382
rect 9884 22260 9940 22270
rect 10220 22260 10276 22316
rect 9884 22258 10276 22260
rect 9884 22206 9886 22258
rect 9938 22206 10276 22258
rect 9884 22204 10276 22206
rect 9884 22194 9940 22204
rect 9548 21810 9716 21812
rect 9548 21758 9550 21810
rect 9602 21758 9716 21810
rect 9548 21756 9716 21758
rect 9772 21924 9828 21934
rect 9548 21746 9604 21756
rect 9772 21586 9828 21868
rect 10220 21924 10276 21934
rect 10332 21924 10388 22988
rect 11452 23042 11508 23054
rect 11452 22990 11454 23042
rect 11506 22990 11508 23042
rect 11340 22932 11396 22942
rect 11228 22372 11284 22382
rect 11228 22278 11284 22316
rect 10276 21868 10388 21924
rect 10444 22148 10500 22158
rect 10444 21924 10500 22092
rect 10892 22148 10948 22158
rect 11340 22148 11396 22876
rect 10892 22054 10948 22092
rect 11228 22092 11396 22148
rect 11452 22482 11508 22990
rect 11452 22430 11454 22482
rect 11506 22430 11508 22482
rect 10220 21858 10276 21868
rect 10444 21858 10500 21868
rect 9772 21534 9774 21586
rect 9826 21534 9828 21586
rect 9772 21522 9828 21534
rect 10108 21698 10164 21710
rect 10108 21646 10110 21698
rect 10162 21646 10164 21698
rect 9660 20804 9716 20814
rect 9548 20692 9604 20702
rect 9324 20690 9604 20692
rect 9324 20638 9550 20690
rect 9602 20638 9604 20690
rect 9324 20636 9604 20638
rect 9212 20244 9268 20636
rect 9212 20188 9492 20244
rect 8652 20020 8708 20030
rect 8540 20018 8708 20020
rect 8540 19966 8654 20018
rect 8706 19966 8708 20018
rect 8540 19964 8708 19966
rect 8428 19926 8484 19964
rect 8540 19460 8596 19470
rect 8540 19366 8596 19404
rect 8316 19294 8318 19346
rect 8370 19294 8372 19346
rect 8316 19282 8372 19294
rect 8652 19012 8708 19964
rect 8876 20018 8932 20030
rect 8876 19966 8878 20018
rect 8930 19966 8932 20018
rect 8764 19906 8820 19918
rect 8764 19854 8766 19906
rect 8818 19854 8820 19906
rect 8764 19348 8820 19854
rect 8876 19458 8932 19966
rect 9436 19908 9492 20188
rect 9548 20132 9604 20636
rect 9660 20242 9716 20748
rect 10108 20804 10164 21646
rect 10444 21700 10500 21710
rect 10444 21698 10724 21700
rect 10444 21646 10446 21698
rect 10498 21646 10724 21698
rect 10444 21644 10724 21646
rect 10444 21634 10500 21644
rect 10556 21476 10612 21486
rect 10108 20738 10164 20748
rect 10220 21474 10612 21476
rect 10220 21422 10558 21474
rect 10610 21422 10612 21474
rect 10220 21420 10612 21422
rect 10220 20692 10276 21420
rect 10556 21410 10612 21420
rect 10668 21140 10724 21644
rect 11004 21474 11060 21486
rect 11004 21422 11006 21474
rect 11058 21422 11060 21474
rect 10668 21084 10948 21140
rect 10220 20690 10388 20692
rect 10220 20638 10222 20690
rect 10274 20638 10388 20690
rect 10220 20636 10388 20638
rect 10220 20626 10276 20636
rect 9660 20190 9662 20242
rect 9714 20190 9716 20242
rect 9660 20178 9716 20190
rect 10220 20356 10276 20366
rect 9548 20066 9604 20076
rect 9772 20130 9828 20142
rect 9772 20078 9774 20130
rect 9826 20078 9828 20130
rect 9548 19908 9604 19918
rect 9436 19906 9604 19908
rect 9436 19854 9550 19906
rect 9602 19854 9604 19906
rect 9436 19852 9604 19854
rect 9548 19842 9604 19852
rect 8876 19406 8878 19458
rect 8930 19406 8932 19458
rect 8876 19394 8932 19406
rect 8764 19282 8820 19292
rect 8764 19012 8820 19022
rect 8652 18956 8764 19012
rect 7980 18674 8372 18676
rect 7980 18622 7982 18674
rect 8034 18622 8372 18674
rect 7980 18620 8372 18622
rect 7980 18610 8036 18620
rect 6972 18470 7028 18508
rect 7532 18564 7588 18574
rect 7532 18470 7588 18508
rect 8316 18562 8372 18620
rect 8764 18674 8820 18956
rect 9324 19012 9380 19022
rect 9324 18918 9380 18956
rect 9772 19010 9828 20078
rect 10220 19796 10276 20300
rect 10332 20244 10388 20636
rect 10332 20150 10388 20188
rect 10444 20690 10500 20702
rect 10444 20638 10446 20690
rect 10498 20638 10500 20690
rect 10444 20020 10500 20638
rect 10332 19796 10388 19806
rect 10220 19794 10388 19796
rect 10220 19742 10334 19794
rect 10386 19742 10388 19794
rect 10220 19740 10388 19742
rect 10332 19730 10388 19740
rect 9772 18958 9774 19010
rect 9826 18958 9828 19010
rect 8764 18622 8766 18674
rect 8818 18622 8820 18674
rect 8764 18610 8820 18622
rect 8316 18510 8318 18562
rect 8370 18510 8372 18562
rect 8316 18498 8372 18510
rect 9772 18564 9828 18958
rect 10220 19012 10276 19022
rect 10220 18918 10276 18956
rect 9772 18498 9828 18508
rect 10220 18788 10276 18798
rect 8540 18450 8596 18462
rect 8540 18398 8542 18450
rect 8594 18398 8596 18450
rect 6972 18228 7028 18238
rect 6748 18226 7028 18228
rect 6748 18174 6974 18226
rect 7026 18174 7028 18226
rect 6748 18172 7028 18174
rect 6972 18162 7028 18172
rect 6524 17778 6692 17780
rect 6524 17726 6526 17778
rect 6578 17726 6692 17778
rect 6524 17724 6692 17726
rect 6524 17714 6580 17724
rect 4732 17666 5124 17668
rect 4732 17614 4734 17666
rect 4786 17614 5124 17666
rect 4732 17612 5124 17614
rect 4732 17602 4788 17612
rect 3724 17462 3780 17500
rect 2604 17444 2660 17454
rect 2604 16884 2660 17388
rect 4060 17444 4116 17454
rect 4060 17350 4116 17388
rect 5068 17444 5124 17612
rect 5068 17378 5124 17388
rect 2940 17108 2996 17118
rect 2940 17014 2996 17052
rect 2156 16828 2324 16884
rect 2156 16658 2212 16670
rect 2156 16606 2158 16658
rect 2210 16606 2212 16658
rect 2156 16212 2212 16606
rect 2156 16146 2212 16156
rect 2044 15986 2100 15998
rect 2044 15934 2046 15986
rect 2098 15934 2100 15986
rect 2044 15540 2100 15934
rect 2044 15474 2100 15484
rect 2268 12964 2324 16828
rect 2604 16818 2660 16828
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 2940 16212 2996 16222
rect 2940 16098 2996 16156
rect 2940 16046 2942 16098
rect 2994 16046 2996 16098
rect 2940 16034 2996 16046
rect 6636 16100 6692 17724
rect 8540 17668 8596 18398
rect 8988 18452 9044 18462
rect 9548 18452 9604 18462
rect 8988 18450 9604 18452
rect 8988 18398 8990 18450
rect 9042 18398 9550 18450
rect 9602 18398 9604 18450
rect 8988 18396 9604 18398
rect 8988 18386 9044 18396
rect 9548 18386 9604 18396
rect 10220 18450 10276 18732
rect 10220 18398 10222 18450
rect 10274 18398 10276 18450
rect 10220 18386 10276 18398
rect 10444 18450 10500 19964
rect 10780 20244 10836 20254
rect 10444 18398 10446 18450
rect 10498 18398 10500 18450
rect 10444 18386 10500 18398
rect 10668 19124 10724 19134
rect 8540 17602 8596 17612
rect 8876 18338 8932 18350
rect 8876 18286 8878 18338
rect 8930 18286 8932 18338
rect 8876 17666 8932 18286
rect 10668 17778 10724 19068
rect 10780 19122 10836 20188
rect 10892 20132 10948 21084
rect 10892 20066 10948 20076
rect 10892 19908 10948 19918
rect 10892 19814 10948 19852
rect 11004 19684 11060 21422
rect 10892 19628 11060 19684
rect 10892 19236 10948 19628
rect 10892 19170 10948 19180
rect 11004 19234 11060 19246
rect 11004 19182 11006 19234
rect 11058 19182 11060 19234
rect 10780 19070 10782 19122
rect 10834 19070 10836 19122
rect 10780 18788 10836 19070
rect 11004 19124 11060 19182
rect 11004 19058 11060 19068
rect 10780 18722 10836 18732
rect 10668 17726 10670 17778
rect 10722 17726 10724 17778
rect 8876 17614 8878 17666
rect 8930 17614 8932 17666
rect 8876 17602 8932 17614
rect 9548 17668 9604 17678
rect 9772 17668 9828 17678
rect 9548 17666 9828 17668
rect 9548 17614 9550 17666
rect 9602 17614 9774 17666
rect 9826 17614 9828 17666
rect 9548 17612 9828 17614
rect 9548 17602 9604 17612
rect 9772 17602 9828 17612
rect 10332 17668 10388 17678
rect 10108 17554 10164 17566
rect 10108 17502 10110 17554
rect 10162 17502 10164 17554
rect 8540 17442 8596 17454
rect 8540 17390 8542 17442
rect 8594 17390 8596 17442
rect 8540 17332 8596 17390
rect 8540 17266 8596 17276
rect 8988 17442 9044 17454
rect 8988 17390 8990 17442
rect 9042 17390 9044 17442
rect 7308 16772 7364 16782
rect 6748 16100 6804 16110
rect 6636 16098 6804 16100
rect 6636 16046 6750 16098
rect 6802 16046 6804 16098
rect 6636 16044 6804 16046
rect 6748 16034 6804 16044
rect 7308 16098 7364 16716
rect 8988 16772 9044 17390
rect 9100 17442 9156 17454
rect 9100 17390 9102 17442
rect 9154 17390 9156 17442
rect 9100 17332 9156 17390
rect 9100 17266 9156 17276
rect 9548 17444 9604 17454
rect 8988 16706 9044 16716
rect 7308 16046 7310 16098
rect 7362 16046 7364 16098
rect 7308 16034 7364 16046
rect 9548 15540 9604 17388
rect 9996 17442 10052 17454
rect 9996 17390 9998 17442
rect 10050 17390 10052 17442
rect 9996 17108 10052 17390
rect 9996 17042 10052 17052
rect 10108 17106 10164 17502
rect 10108 17054 10110 17106
rect 10162 17054 10164 17106
rect 10108 16996 10164 17054
rect 10108 16930 10164 16940
rect 10332 16994 10388 17612
rect 10668 17668 10724 17726
rect 10668 17602 10724 17612
rect 10780 18452 10836 18462
rect 11116 18452 11172 18462
rect 10780 17666 10836 18396
rect 10780 17614 10782 17666
rect 10834 17614 10836 17666
rect 10332 16942 10334 16994
rect 10386 16942 10388 16994
rect 10332 16930 10388 16942
rect 10444 17108 10500 17118
rect 10332 16324 10388 16334
rect 10444 16324 10500 17052
rect 10780 17108 10836 17614
rect 10780 17042 10836 17052
rect 10892 18450 11172 18452
rect 10892 18398 11118 18450
rect 11170 18398 11172 18450
rect 10892 18396 11172 18398
rect 10892 16660 10948 18396
rect 11116 18386 11172 18396
rect 11116 18226 11172 18238
rect 11116 18174 11118 18226
rect 11170 18174 11172 18226
rect 11004 17780 11060 17790
rect 11004 16882 11060 17724
rect 11004 16830 11006 16882
rect 11058 16830 11060 16882
rect 11004 16818 11060 16830
rect 11116 16770 11172 18174
rect 11116 16718 11118 16770
rect 11170 16718 11172 16770
rect 11116 16706 11172 16718
rect 10892 16594 10948 16604
rect 11228 16548 11284 22092
rect 11340 21924 11396 21934
rect 11340 18228 11396 21868
rect 11452 21700 11508 22430
rect 12908 22484 12964 22494
rect 12012 22370 12068 22382
rect 12012 22318 12014 22370
rect 12066 22318 12068 22370
rect 11900 22260 11956 22270
rect 11900 22146 11956 22204
rect 11900 22094 11902 22146
rect 11954 22094 11956 22146
rect 11900 22082 11956 22094
rect 11452 21634 11508 21644
rect 11788 21028 11844 21038
rect 12012 21028 12068 22318
rect 12684 22372 12740 22382
rect 12572 21700 12628 21710
rect 12572 21606 12628 21644
rect 12348 21586 12404 21598
rect 12348 21534 12350 21586
rect 12402 21534 12404 21586
rect 12348 21028 12404 21534
rect 11788 21026 12404 21028
rect 11788 20974 11790 21026
rect 11842 20974 12404 21026
rect 11788 20972 12404 20974
rect 12684 21026 12740 22316
rect 12908 22258 12964 22428
rect 12908 22206 12910 22258
rect 12962 22206 12964 22258
rect 12908 22194 12964 22206
rect 13692 22484 13748 22494
rect 13468 22148 13524 22158
rect 12908 21812 12964 21822
rect 12908 21718 12964 21756
rect 13468 21586 13524 22092
rect 13468 21534 13470 21586
rect 13522 21534 13524 21586
rect 13468 21522 13524 21534
rect 13692 21810 13748 22428
rect 14140 22372 14196 28140
rect 14364 25506 14420 28588
rect 15148 28644 15204 28654
rect 15148 28550 15204 28588
rect 15932 28642 15988 34972
rect 16268 35026 16324 35646
rect 16492 35700 16548 35710
rect 16492 35364 16548 35644
rect 16492 35298 16548 35308
rect 16268 34974 16270 35026
rect 16322 34974 16324 35026
rect 16268 34962 16324 34974
rect 16380 35252 16436 35262
rect 16380 35028 16436 35196
rect 16044 34916 16100 34926
rect 16044 34822 16100 34860
rect 16268 34804 16324 34814
rect 16268 34690 16324 34748
rect 16268 34638 16270 34690
rect 16322 34638 16324 34690
rect 16268 34244 16324 34638
rect 16380 34692 16436 34972
rect 16492 34916 16548 34926
rect 16492 34822 16548 34860
rect 16716 34692 16772 36204
rect 17164 35924 17220 37774
rect 17388 37492 17444 37502
rect 17388 37398 17444 37436
rect 16828 35868 17220 35924
rect 16828 35700 16884 35868
rect 16828 35634 16884 35644
rect 16940 35700 16996 35710
rect 17500 35700 17556 37998
rect 18060 37268 18116 37278
rect 17948 37266 18116 37268
rect 17948 37214 18062 37266
rect 18114 37214 18116 37266
rect 17948 37212 18116 37214
rect 17836 35700 17892 35710
rect 16940 35698 17332 35700
rect 16940 35646 16942 35698
rect 16994 35646 17332 35698
rect 16940 35644 17332 35646
rect 17500 35644 17836 35700
rect 16940 35634 16996 35644
rect 17164 35476 17220 35486
rect 16828 34916 16884 34926
rect 16828 34822 16884 34860
rect 16380 34626 16436 34636
rect 16492 34636 16772 34692
rect 16156 34188 16324 34244
rect 16156 32452 16212 34188
rect 16268 34018 16324 34030
rect 16268 33966 16270 34018
rect 16322 33966 16324 34018
rect 16268 33348 16324 33966
rect 16492 33458 16548 34636
rect 16940 34356 16996 34366
rect 16940 34262 16996 34300
rect 16716 34242 16772 34254
rect 16716 34190 16718 34242
rect 16770 34190 16772 34242
rect 16604 34130 16660 34142
rect 16604 34078 16606 34130
rect 16658 34078 16660 34130
rect 16604 34020 16660 34078
rect 16604 33572 16660 33964
rect 16604 33506 16660 33516
rect 16492 33406 16494 33458
rect 16546 33406 16548 33458
rect 16492 33394 16548 33406
rect 16380 33348 16436 33358
rect 16268 33346 16436 33348
rect 16268 33294 16382 33346
rect 16434 33294 16436 33346
rect 16268 33292 16436 33294
rect 16380 33282 16436 33292
rect 16604 33348 16660 33358
rect 16604 32788 16660 33292
rect 16716 33236 16772 34190
rect 17052 33460 17108 33470
rect 17052 33346 17108 33404
rect 17052 33294 17054 33346
rect 17106 33294 17108 33346
rect 17052 33282 17108 33294
rect 16716 33170 16772 33180
rect 16828 32788 16884 32798
rect 16492 32786 16884 32788
rect 16492 32734 16830 32786
rect 16882 32734 16884 32786
rect 16492 32732 16884 32734
rect 16380 32452 16436 32462
rect 16156 32450 16436 32452
rect 16156 32398 16382 32450
rect 16434 32398 16436 32450
rect 16156 32396 16436 32398
rect 16156 30100 16212 30110
rect 16156 30006 16212 30044
rect 16156 29428 16212 29438
rect 16156 29334 16212 29372
rect 16268 29316 16324 32396
rect 16380 32386 16436 32396
rect 16492 30324 16548 32732
rect 16828 32722 16884 32732
rect 17164 31892 17220 35420
rect 17276 35252 17332 35644
rect 17836 35606 17892 35644
rect 17388 35588 17444 35598
rect 17388 35494 17444 35532
rect 17948 35588 18004 37212
rect 18060 37202 18116 37212
rect 18060 36148 18116 36158
rect 18116 36092 18228 36148
rect 18060 36082 18116 36092
rect 17948 35522 18004 35532
rect 18172 35586 18228 36092
rect 18284 35924 18340 38612
rect 18732 38612 18900 38668
rect 18732 38164 18788 38612
rect 19516 38276 19572 41200
rect 19516 38210 19572 38220
rect 20188 38274 20244 41200
rect 20860 39620 20916 41200
rect 20860 39564 21364 39620
rect 20188 38222 20190 38274
rect 20242 38222 20244 38274
rect 20188 38210 20244 38222
rect 18732 38162 19012 38164
rect 18732 38110 18734 38162
rect 18786 38110 19012 38162
rect 18732 38108 19012 38110
rect 18732 38098 18788 38108
rect 18956 37490 19012 38108
rect 21308 38162 21364 39564
rect 21532 38668 21588 41200
rect 21532 38612 21700 38668
rect 21308 38110 21310 38162
rect 21362 38110 21364 38162
rect 21308 38098 21364 38110
rect 18956 37438 18958 37490
rect 19010 37438 19012 37490
rect 18956 37426 19012 37438
rect 19068 37996 19460 38052
rect 18620 37154 18676 37166
rect 18620 37102 18622 37154
rect 18674 37102 18676 37154
rect 18620 36372 18676 37102
rect 18620 36036 18676 36316
rect 18620 35970 18676 35980
rect 18284 35858 18340 35868
rect 18172 35534 18174 35586
rect 18226 35534 18228 35586
rect 17276 35196 18116 35252
rect 17500 34916 17556 34926
rect 17556 34860 17668 34916
rect 17500 34822 17556 34860
rect 17500 34354 17556 34366
rect 17500 34302 17502 34354
rect 17554 34302 17556 34354
rect 17388 34244 17444 34254
rect 17388 34130 17444 34188
rect 17388 34078 17390 34130
rect 17442 34078 17444 34130
rect 17388 34066 17444 34078
rect 17500 33348 17556 34302
rect 17612 34130 17668 34860
rect 17724 34914 17780 34926
rect 17724 34862 17726 34914
rect 17778 34862 17780 34914
rect 17724 34356 17780 34862
rect 18060 34914 18116 35196
rect 18060 34862 18062 34914
rect 18114 34862 18116 34914
rect 18060 34850 18116 34862
rect 18172 34916 18228 35534
rect 18172 34850 18228 34860
rect 18284 35700 18340 35710
rect 18284 34802 18340 35644
rect 18732 35588 18788 35598
rect 18508 35586 18788 35588
rect 18508 35534 18734 35586
rect 18786 35534 18788 35586
rect 18508 35532 18788 35534
rect 18396 35140 18452 35150
rect 18396 34914 18452 35084
rect 18396 34862 18398 34914
rect 18450 34862 18452 34914
rect 18396 34850 18452 34862
rect 18284 34750 18286 34802
rect 18338 34750 18340 34802
rect 18284 34738 18340 34750
rect 18508 34580 18564 35532
rect 18732 35522 18788 35532
rect 18844 35028 18900 35038
rect 18732 34916 18788 34926
rect 18620 34692 18676 34702
rect 18620 34598 18676 34636
rect 17724 34290 17780 34300
rect 18396 34524 18564 34580
rect 17612 34078 17614 34130
rect 17666 34078 17668 34130
rect 17612 34066 17668 34078
rect 17836 33572 17892 33582
rect 17612 33348 17668 33358
rect 17500 33346 17668 33348
rect 17500 33294 17614 33346
rect 17666 33294 17668 33346
rect 17500 33292 17668 33294
rect 17612 32564 17668 33292
rect 17836 33234 17892 33516
rect 18396 33460 18452 34524
rect 18508 34356 18564 34366
rect 18508 34262 18564 34300
rect 18732 34354 18788 34860
rect 18844 34802 18900 34972
rect 18844 34750 18846 34802
rect 18898 34750 18900 34802
rect 18844 34738 18900 34750
rect 18956 34802 19012 34814
rect 18956 34750 18958 34802
rect 19010 34750 19012 34802
rect 18956 34580 19012 34750
rect 18732 34302 18734 34354
rect 18786 34302 18788 34354
rect 18732 34290 18788 34302
rect 18844 34524 19012 34580
rect 18844 34244 18900 34524
rect 19068 34356 19124 37996
rect 19180 37828 19236 37838
rect 19180 37826 19348 37828
rect 19180 37774 19182 37826
rect 19234 37774 19348 37826
rect 19180 37772 19348 37774
rect 19180 37762 19236 37772
rect 19292 37604 19348 37772
rect 19404 37826 19460 37996
rect 19404 37774 19406 37826
rect 19458 37774 19460 37826
rect 19404 37762 19460 37774
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19292 37548 19572 37604
rect 19836 37594 20100 37604
rect 19292 37380 19348 37390
rect 19292 37378 19460 37380
rect 19292 37326 19294 37378
rect 19346 37326 19460 37378
rect 19292 37324 19460 37326
rect 19292 37314 19348 37324
rect 19180 35924 19236 35934
rect 19180 35700 19236 35868
rect 19404 35812 19460 37324
rect 19516 37268 19572 37548
rect 19516 37174 19572 37212
rect 20188 37268 20244 37278
rect 20188 37266 21476 37268
rect 20188 37214 20190 37266
rect 20242 37214 21476 37266
rect 20188 37212 21476 37214
rect 20188 37202 20244 37212
rect 21420 36594 21476 37212
rect 21420 36542 21422 36594
rect 21474 36542 21476 36594
rect 21420 36530 21476 36542
rect 20524 36372 20580 36382
rect 20524 36278 20580 36316
rect 19628 36260 19684 36270
rect 19628 36166 19684 36204
rect 20188 36258 20244 36270
rect 20188 36206 20190 36258
rect 20242 36206 20244 36258
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19628 35812 19684 35822
rect 19404 35756 19572 35812
rect 19180 35698 19460 35700
rect 19180 35646 19182 35698
rect 19234 35646 19460 35698
rect 19180 35644 19460 35646
rect 19180 35634 19236 35644
rect 19180 35140 19236 35150
rect 19236 35084 19348 35140
rect 19180 35074 19236 35084
rect 18844 34178 18900 34188
rect 18956 34300 19124 34356
rect 18620 34018 18676 34030
rect 18620 33966 18622 34018
rect 18674 33966 18676 34018
rect 18620 33572 18676 33966
rect 18620 33516 18900 33572
rect 18396 33404 18676 33460
rect 17836 33182 17838 33234
rect 17890 33182 17892 33234
rect 17724 32564 17780 32574
rect 17612 32562 17780 32564
rect 17612 32510 17726 32562
rect 17778 32510 17780 32562
rect 17612 32508 17780 32510
rect 17724 32498 17780 32508
rect 17836 32564 17892 33182
rect 18396 33236 18452 33246
rect 17836 32498 17892 32508
rect 18284 32674 18340 32686
rect 18284 32622 18286 32674
rect 18338 32622 18340 32674
rect 16940 31836 17220 31892
rect 16828 31668 16884 31678
rect 16716 31220 16772 31230
rect 16716 31126 16772 31164
rect 16604 31106 16660 31118
rect 16604 31054 16606 31106
rect 16658 31054 16660 31106
rect 16604 30884 16660 31054
rect 16828 31106 16884 31612
rect 16828 31054 16830 31106
rect 16882 31054 16884 31106
rect 16828 31042 16884 31054
rect 16604 30818 16660 30828
rect 16940 30324 16996 31836
rect 17276 31780 17332 31790
rect 17276 31686 17332 31724
rect 16492 30268 16772 30324
rect 16380 29652 16436 29662
rect 16380 29426 16436 29596
rect 16380 29374 16382 29426
rect 16434 29374 16436 29426
rect 16380 29362 16436 29374
rect 16268 29250 16324 29260
rect 16716 28868 16772 30268
rect 16716 28774 16772 28812
rect 16828 30268 16996 30324
rect 17052 31666 17108 31678
rect 17052 31614 17054 31666
rect 17106 31614 17108 31666
rect 16828 29428 16884 30268
rect 15932 28590 15934 28642
rect 15986 28590 15988 28642
rect 14700 28082 14756 28094
rect 14700 28030 14702 28082
rect 14754 28030 14756 28082
rect 14700 25730 14756 28030
rect 15932 28084 15988 28590
rect 16828 28756 16884 29372
rect 16268 28532 16324 28542
rect 16268 28438 16324 28476
rect 15932 28018 15988 28028
rect 16604 28084 16660 28094
rect 16604 27990 16660 28028
rect 15932 27748 15988 27758
rect 15988 27692 16436 27748
rect 15932 27654 15988 27692
rect 14700 25678 14702 25730
rect 14754 25678 14756 25730
rect 14700 25666 14756 25678
rect 14812 27636 14868 27646
rect 14812 25844 14868 27580
rect 15372 27634 15428 27646
rect 15372 27582 15374 27634
rect 15426 27582 15428 27634
rect 15260 26292 15316 26302
rect 15260 25844 15316 26236
rect 14812 25788 15316 25844
rect 14812 25618 14868 25788
rect 14812 25566 14814 25618
rect 14866 25566 14868 25618
rect 14812 25554 14868 25566
rect 14924 25620 14980 25630
rect 14364 25454 14366 25506
rect 14418 25454 14420 25506
rect 14364 25442 14420 25454
rect 14924 24722 14980 25564
rect 15260 25618 15316 25788
rect 15260 25566 15262 25618
rect 15314 25566 15316 25618
rect 15260 25554 15316 25566
rect 15372 25620 15428 27582
rect 16268 26852 16324 26862
rect 16044 26850 16324 26852
rect 16044 26798 16270 26850
rect 16322 26798 16324 26850
rect 16044 26796 16324 26798
rect 16044 26514 16100 26796
rect 16268 26786 16324 26796
rect 16044 26462 16046 26514
rect 16098 26462 16100 26514
rect 16044 26450 16100 26462
rect 15372 25554 15428 25564
rect 15484 26290 15540 26302
rect 15484 26238 15486 26290
rect 15538 26238 15540 26290
rect 15484 25284 15540 26238
rect 15932 26292 15988 26302
rect 15932 26198 15988 26236
rect 15820 25732 15876 25742
rect 15708 25284 15764 25294
rect 15484 25228 15708 25284
rect 15708 25190 15764 25228
rect 15820 25172 15876 25676
rect 16380 25620 16436 27692
rect 16828 27300 16884 28700
rect 16940 30100 16996 30110
rect 16940 28754 16996 30044
rect 17052 29876 17108 31614
rect 18284 31220 18340 32622
rect 18396 32676 18452 33180
rect 18396 32610 18452 32620
rect 18620 31778 18676 33404
rect 18844 33346 18900 33516
rect 18844 33294 18846 33346
rect 18898 33294 18900 33346
rect 18844 33282 18900 33294
rect 18732 33234 18788 33246
rect 18732 33182 18734 33234
rect 18786 33182 18788 33234
rect 18732 33124 18788 33182
rect 18844 33124 18900 33134
rect 18732 33068 18844 33124
rect 18620 31726 18622 31778
rect 18674 31726 18676 31778
rect 18396 31668 18452 31678
rect 18396 31574 18452 31612
rect 18284 31154 18340 31164
rect 18508 31108 18564 31118
rect 18508 31014 18564 31052
rect 17500 30996 17556 31006
rect 17500 30902 17556 30940
rect 17948 30996 18004 31006
rect 18172 30996 18228 31006
rect 17948 30994 18116 30996
rect 17948 30942 17950 30994
rect 18002 30942 18116 30994
rect 17948 30940 18116 30942
rect 17948 30930 18004 30940
rect 17052 29810 17108 29820
rect 17164 30884 17220 30894
rect 17164 30212 17220 30828
rect 17724 30882 17780 30894
rect 17724 30830 17726 30882
rect 17778 30830 17780 30882
rect 17388 30324 17444 30334
rect 17388 30230 17444 30268
rect 17164 29652 17220 30156
rect 17612 30098 17668 30110
rect 17612 30046 17614 30098
rect 17666 30046 17668 30098
rect 17612 29876 17668 30046
rect 17724 30100 17780 30830
rect 18060 30884 18116 30940
rect 17948 30212 18004 30222
rect 17724 30034 17780 30044
rect 17836 30210 18004 30212
rect 17836 30158 17950 30210
rect 18002 30158 18004 30210
rect 17836 30156 18004 30158
rect 17612 29810 17668 29820
rect 17612 29652 17668 29662
rect 17836 29652 17892 30156
rect 17948 30146 18004 30156
rect 17220 29596 17556 29652
rect 17164 29558 17220 29596
rect 17500 29538 17556 29596
rect 17612 29650 17892 29652
rect 17612 29598 17614 29650
rect 17666 29598 17892 29650
rect 17612 29596 17892 29598
rect 17612 29586 17668 29596
rect 17500 29486 17502 29538
rect 17554 29486 17556 29538
rect 17500 29474 17556 29486
rect 16940 28702 16942 28754
rect 16994 28702 16996 28754
rect 16940 28690 16996 28702
rect 17388 29428 17444 29438
rect 17388 28642 17444 29372
rect 17612 29428 17668 29438
rect 17612 29202 17668 29372
rect 17612 29150 17614 29202
rect 17666 29150 17668 29202
rect 17612 29138 17668 29150
rect 17388 28590 17390 28642
rect 17442 28590 17444 28642
rect 17388 28578 17444 28590
rect 17724 28868 17780 28878
rect 17276 28532 17332 28542
rect 17276 28438 17332 28476
rect 17164 28420 17220 28430
rect 17052 27300 17108 27310
rect 16828 27298 17108 27300
rect 16828 27246 17054 27298
rect 17106 27246 17108 27298
rect 16828 27244 17108 27246
rect 17052 27234 17108 27244
rect 16940 26964 16996 26974
rect 16492 26292 16548 26302
rect 16492 26198 16548 26236
rect 16380 25618 16660 25620
rect 16380 25566 16382 25618
rect 16434 25566 16660 25618
rect 16380 25564 16660 25566
rect 16380 25554 16436 25564
rect 16604 25506 16660 25564
rect 16604 25454 16606 25506
rect 16658 25454 16660 25506
rect 16604 25442 16660 25454
rect 15820 24946 15876 25116
rect 15820 24894 15822 24946
rect 15874 24894 15876 24946
rect 15820 24882 15876 24894
rect 14924 24670 14926 24722
rect 14978 24670 14980 24722
rect 14924 24658 14980 24670
rect 15260 24834 15316 24846
rect 15260 24782 15262 24834
rect 15314 24782 15316 24834
rect 14476 24052 14532 24062
rect 14532 23996 14756 24052
rect 14476 23958 14532 23996
rect 14700 23938 14756 23996
rect 14700 23886 14702 23938
rect 14754 23886 14756 23938
rect 14700 23874 14756 23886
rect 13692 21758 13694 21810
rect 13746 21758 13748 21810
rect 12684 20974 12686 21026
rect 12738 20974 12740 21026
rect 11788 20962 11844 20972
rect 12684 20962 12740 20974
rect 13468 21364 13524 21374
rect 12124 20802 12180 20814
rect 12124 20750 12126 20802
rect 12178 20750 12180 20802
rect 11676 20692 11732 20702
rect 11564 20690 11732 20692
rect 11564 20638 11678 20690
rect 11730 20638 11732 20690
rect 11564 20636 11732 20638
rect 11564 19346 11620 20636
rect 11676 20626 11732 20636
rect 11564 19294 11566 19346
rect 11618 19294 11620 19346
rect 11564 19282 11620 19294
rect 11676 19234 11732 19246
rect 11676 19182 11678 19234
rect 11730 19182 11732 19234
rect 11452 19122 11508 19134
rect 11452 19070 11454 19122
rect 11506 19070 11508 19122
rect 11452 18452 11508 19070
rect 11676 18788 11732 19182
rect 11676 18722 11732 18732
rect 11900 19234 11956 19246
rect 11900 19182 11902 19234
rect 11954 19182 11956 19234
rect 11452 18386 11508 18396
rect 11340 18162 11396 18172
rect 11452 18226 11508 18238
rect 11788 18228 11844 18238
rect 11452 18174 11454 18226
rect 11506 18174 11508 18226
rect 11452 18004 11508 18174
rect 11452 17938 11508 17948
rect 11564 18226 11844 18228
rect 11564 18174 11790 18226
rect 11842 18174 11844 18226
rect 11564 18172 11844 18174
rect 11452 17780 11508 17790
rect 11564 17780 11620 18172
rect 11788 18162 11844 18172
rect 11508 17724 11620 17780
rect 11900 17778 11956 19182
rect 12124 19234 12180 20750
rect 12348 20804 12404 20814
rect 12348 20710 12404 20748
rect 13468 20804 13524 21308
rect 13468 20710 13524 20748
rect 13692 20802 13748 21758
rect 14028 22316 14196 22372
rect 15148 23716 15204 23726
rect 15260 23716 15316 24782
rect 16380 24724 16436 24734
rect 16380 24610 16436 24668
rect 16380 24558 16382 24610
rect 16434 24558 16436 24610
rect 15204 23660 15316 23716
rect 15372 23938 15428 23950
rect 15372 23886 15374 23938
rect 15426 23886 15428 23938
rect 14028 21812 14084 22316
rect 14140 22148 14196 22158
rect 14588 22148 14644 22158
rect 14140 22146 14644 22148
rect 14140 22094 14142 22146
rect 14194 22094 14590 22146
rect 14642 22094 14644 22146
rect 14140 22092 14644 22094
rect 14140 22082 14196 22092
rect 14028 21746 14084 21756
rect 14476 21698 14532 22092
rect 14588 22082 14644 22092
rect 14700 22148 14756 22158
rect 14700 21810 14756 22092
rect 14700 21758 14702 21810
rect 14754 21758 14756 21810
rect 14700 21746 14756 21758
rect 14476 21646 14478 21698
rect 14530 21646 14532 21698
rect 14364 21588 14420 21598
rect 14252 21586 14420 21588
rect 14252 21534 14366 21586
rect 14418 21534 14420 21586
rect 14252 21532 14420 21534
rect 13692 20750 13694 20802
rect 13746 20750 13748 20802
rect 13692 20738 13748 20750
rect 13916 20802 13972 20814
rect 13916 20750 13918 20802
rect 13970 20750 13972 20802
rect 13580 20580 13636 20590
rect 13468 20578 13636 20580
rect 13468 20526 13582 20578
rect 13634 20526 13636 20578
rect 13468 20524 13636 20526
rect 12236 19908 12292 19918
rect 12684 19908 12740 19918
rect 12236 19906 12740 19908
rect 12236 19854 12238 19906
rect 12290 19854 12686 19906
rect 12738 19854 12740 19906
rect 12236 19852 12740 19854
rect 12236 19684 12292 19852
rect 12236 19618 12292 19628
rect 12124 19182 12126 19234
rect 12178 19182 12180 19234
rect 12012 18562 12068 18574
rect 12012 18510 12014 18562
rect 12066 18510 12068 18562
rect 12012 18452 12068 18510
rect 12012 18386 12068 18396
rect 12124 18338 12180 19182
rect 12460 19348 12516 19358
rect 12460 19234 12516 19292
rect 12460 19182 12462 19234
rect 12514 19182 12516 19234
rect 12460 19170 12516 19182
rect 12684 19124 12740 19852
rect 12796 19460 12852 19470
rect 12796 19458 13188 19460
rect 12796 19406 12798 19458
rect 12850 19406 13188 19458
rect 12796 19404 13188 19406
rect 12796 19394 12852 19404
rect 12908 19236 12964 19246
rect 12908 19142 12964 19180
rect 12684 19058 12740 19068
rect 12796 19010 12852 19022
rect 12796 18958 12798 19010
rect 12850 18958 12852 19010
rect 12796 18452 12852 18958
rect 12684 18396 12796 18452
rect 12124 18286 12126 18338
rect 12178 18286 12180 18338
rect 12124 18274 12180 18286
rect 12572 18340 12628 18350
rect 12572 18246 12628 18284
rect 12460 18228 12516 18238
rect 12348 18226 12516 18228
rect 12348 18174 12462 18226
rect 12514 18174 12516 18226
rect 12348 18172 12516 18174
rect 11900 17726 11902 17778
rect 11954 17726 11956 17778
rect 11452 17686 11508 17724
rect 11900 17714 11956 17726
rect 12236 18116 12292 18126
rect 11788 17668 11844 17678
rect 11788 17574 11844 17612
rect 12124 17666 12180 17678
rect 12124 17614 12126 17666
rect 12178 17614 12180 17666
rect 12124 17444 12180 17614
rect 12236 17666 12292 18060
rect 12236 17614 12238 17666
rect 12290 17614 12292 17666
rect 12236 17602 12292 17614
rect 12348 17444 12404 18172
rect 12460 18162 12516 18172
rect 12124 17388 12404 17444
rect 12572 17666 12628 17678
rect 12572 17614 12574 17666
rect 12626 17614 12628 17666
rect 12012 17332 12068 17342
rect 11900 17108 11956 17118
rect 11788 17052 11900 17108
rect 11788 16994 11844 17052
rect 11900 17042 11956 17052
rect 12012 17108 12068 17276
rect 12012 17106 12292 17108
rect 12012 17054 12014 17106
rect 12066 17054 12292 17106
rect 12012 17052 12292 17054
rect 12012 17042 12068 17052
rect 11788 16942 11790 16994
rect 11842 16942 11844 16994
rect 11788 16930 11844 16942
rect 11228 16482 11284 16492
rect 11900 16770 11956 16782
rect 11900 16718 11902 16770
rect 11954 16718 11956 16770
rect 10332 16322 10500 16324
rect 10332 16270 10334 16322
rect 10386 16270 10500 16322
rect 10332 16268 10500 16270
rect 10332 16258 10388 16268
rect 11116 15988 11172 15998
rect 9548 15426 9604 15484
rect 9660 15874 9716 15886
rect 9660 15822 9662 15874
rect 9714 15822 9716 15874
rect 9660 15538 9716 15822
rect 10668 15874 10724 15886
rect 10668 15822 10670 15874
rect 10722 15822 10724 15874
rect 9660 15486 9662 15538
rect 9714 15486 9716 15538
rect 9660 15474 9716 15486
rect 10108 15540 10164 15550
rect 10108 15446 10164 15484
rect 9548 15374 9550 15426
rect 9602 15374 9604 15426
rect 9548 15362 9604 15374
rect 10668 15314 10724 15822
rect 10668 15262 10670 15314
rect 10722 15262 10724 15314
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 10108 14532 10164 14542
rect 9996 14476 10108 14532
rect 7532 14420 7588 14430
rect 7532 14326 7588 14364
rect 8428 14420 8484 14430
rect 8428 14326 8484 14364
rect 7196 14308 7252 14318
rect 7420 14308 7476 14318
rect 2940 13860 2996 13870
rect 2940 13074 2996 13804
rect 5068 13860 5124 13870
rect 5068 13766 5124 13804
rect 5404 13748 5460 13758
rect 5404 13746 5684 13748
rect 5404 13694 5406 13746
rect 5458 13694 5684 13746
rect 5404 13692 5684 13694
rect 5404 13682 5460 13692
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 2940 13022 2942 13074
rect 2994 13022 2996 13074
rect 2940 13010 2996 13022
rect 5068 13188 5124 13198
rect 5068 13074 5124 13132
rect 5068 13022 5070 13074
rect 5122 13022 5124 13074
rect 5068 13010 5124 13022
rect 5628 13074 5684 13692
rect 6076 13636 6132 13646
rect 6076 13542 6132 13580
rect 7196 13636 7252 14252
rect 5628 13022 5630 13074
rect 5682 13022 5684 13074
rect 5628 13010 5684 13022
rect 6524 13188 6580 13198
rect 6524 13074 6580 13132
rect 7196 13186 7252 13580
rect 7196 13134 7198 13186
rect 7250 13134 7252 13186
rect 7196 13122 7252 13134
rect 7308 14306 7476 14308
rect 7308 14254 7422 14306
rect 7474 14254 7476 14306
rect 7308 14252 7476 14254
rect 7308 13188 7364 14252
rect 7420 14242 7476 14252
rect 7644 14306 7700 14318
rect 7644 14254 7646 14306
rect 7698 14254 7700 14306
rect 7532 13188 7588 13198
rect 7644 13188 7700 14254
rect 7868 14308 7924 14318
rect 8316 14308 8372 14318
rect 7868 14214 7924 14252
rect 8204 14306 8372 14308
rect 8204 14254 8318 14306
rect 8370 14254 8372 14306
rect 8204 14252 8372 14254
rect 8204 13858 8260 14252
rect 8316 14242 8372 14252
rect 8204 13806 8206 13858
rect 8258 13806 8260 13858
rect 8204 13794 8260 13806
rect 8988 13748 9044 13758
rect 8988 13654 9044 13692
rect 9660 13748 9716 13758
rect 9660 13636 9716 13692
rect 9996 13636 10052 14476
rect 10108 14466 10164 14476
rect 10668 14532 10724 15262
rect 11116 15314 11172 15932
rect 11900 15988 11956 16718
rect 12236 16210 12292 17052
rect 12460 16884 12516 16894
rect 12460 16790 12516 16828
rect 12460 16660 12516 16670
rect 12460 16322 12516 16604
rect 12460 16270 12462 16322
rect 12514 16270 12516 16322
rect 12460 16258 12516 16270
rect 12572 16324 12628 17614
rect 12684 17556 12740 18396
rect 12796 18386 12852 18396
rect 12908 18900 12964 18910
rect 12684 16994 12740 17500
rect 12684 16942 12686 16994
rect 12738 16942 12740 16994
rect 12684 16930 12740 16942
rect 12796 18116 12852 18126
rect 12908 18116 12964 18844
rect 13132 18674 13188 19404
rect 13468 19236 13524 20524
rect 13580 20514 13636 20524
rect 13916 19348 13972 20750
rect 14252 20692 14308 21532
rect 14364 21522 14420 21532
rect 14476 21252 14532 21646
rect 14924 21364 14980 21374
rect 14924 21270 14980 21308
rect 14028 20244 14084 20254
rect 14028 19908 14084 20188
rect 14140 20132 14196 20142
rect 14252 20132 14308 20636
rect 14364 21196 14532 21252
rect 14364 20690 14420 21196
rect 14476 21028 14532 21038
rect 14476 20934 14532 20972
rect 14364 20638 14366 20690
rect 14418 20638 14420 20690
rect 14364 20580 14420 20638
rect 14364 20524 14644 20580
rect 14140 20130 14532 20132
rect 14140 20078 14142 20130
rect 14194 20078 14532 20130
rect 14140 20076 14532 20078
rect 14140 20066 14196 20076
rect 14028 19852 14196 19908
rect 13916 19282 13972 19292
rect 13132 18622 13134 18674
rect 13186 18622 13188 18674
rect 13132 18610 13188 18622
rect 13356 18788 13412 18798
rect 13356 18674 13412 18732
rect 13356 18622 13358 18674
rect 13410 18622 13412 18674
rect 13356 18610 13412 18622
rect 12852 18060 12964 18116
rect 13020 18450 13076 18462
rect 13020 18398 13022 18450
rect 13074 18398 13076 18450
rect 12236 16158 12238 16210
rect 12290 16158 12292 16210
rect 12236 16146 12292 16158
rect 11900 15922 11956 15932
rect 12572 15986 12628 16268
rect 12796 16882 12852 18060
rect 13020 17892 13076 18398
rect 13020 17826 13076 17836
rect 13244 18338 13300 18350
rect 13244 18286 13246 18338
rect 13298 18286 13300 18338
rect 13244 17108 13300 18286
rect 13468 18228 13524 19180
rect 13692 19122 13748 19134
rect 13692 19070 13694 19122
rect 13746 19070 13748 19122
rect 13692 18900 13748 19070
rect 13916 19124 13972 19134
rect 13916 19030 13972 19068
rect 14028 19122 14084 19134
rect 14028 19070 14030 19122
rect 14082 19070 14084 19122
rect 13692 18834 13748 18844
rect 14028 18788 14084 19070
rect 14028 18722 14084 18732
rect 14028 18562 14084 18574
rect 14028 18510 14030 18562
rect 14082 18510 14084 18562
rect 13580 18450 13636 18462
rect 13580 18398 13582 18450
rect 13634 18398 13636 18450
rect 13580 18340 13636 18398
rect 13916 18340 13972 18350
rect 13580 18338 13972 18340
rect 13580 18286 13918 18338
rect 13970 18286 13972 18338
rect 13580 18284 13972 18286
rect 13916 18274 13972 18284
rect 13468 18172 13860 18228
rect 13468 18004 13524 18014
rect 13468 17890 13524 17948
rect 13468 17838 13470 17890
rect 13522 17838 13524 17890
rect 13468 17780 13524 17838
rect 13804 17890 13860 18172
rect 13804 17838 13806 17890
rect 13858 17838 13860 17890
rect 13804 17826 13860 17838
rect 13468 17714 13524 17724
rect 13468 17556 13524 17566
rect 13524 17500 13636 17556
rect 13468 17490 13524 17500
rect 13580 17442 13636 17500
rect 13580 17390 13582 17442
rect 13634 17390 13636 17442
rect 13580 17378 13636 17390
rect 14028 17444 14084 18510
rect 14140 18564 14196 19852
rect 14252 19796 14308 19806
rect 14252 19458 14308 19740
rect 14252 19406 14254 19458
rect 14306 19406 14308 19458
rect 14252 19394 14308 19406
rect 14476 19458 14532 20076
rect 14476 19406 14478 19458
rect 14530 19406 14532 19458
rect 14476 19394 14532 19406
rect 14588 20020 14644 20524
rect 14588 19124 14644 19964
rect 14588 19058 14644 19068
rect 14700 20018 14756 20030
rect 14700 19966 14702 20018
rect 14754 19966 14756 20018
rect 14700 18900 14756 19966
rect 15036 20018 15092 20030
rect 15036 19966 15038 20018
rect 15090 19966 15092 20018
rect 15036 19796 15092 19966
rect 14700 18834 14756 18844
rect 14924 19740 15036 19796
rect 14252 18564 14308 18574
rect 14140 18562 14308 18564
rect 14140 18510 14254 18562
rect 14306 18510 14308 18562
rect 14140 18508 14308 18510
rect 14252 18498 14308 18508
rect 14924 18562 14980 19740
rect 15036 19730 15092 19740
rect 15148 19684 15204 23660
rect 15372 23156 15428 23886
rect 16380 23604 16436 24558
rect 16380 23538 16436 23548
rect 16828 24612 16884 24622
rect 16268 23380 16324 23390
rect 15372 23090 15428 23100
rect 15932 23378 16324 23380
rect 15932 23326 16270 23378
rect 16322 23326 16324 23378
rect 15932 23324 16324 23326
rect 15932 22484 15988 23324
rect 16268 23314 16324 23324
rect 16828 23380 16884 24556
rect 16156 23154 16212 23166
rect 16156 23102 16158 23154
rect 16210 23102 16212 23154
rect 16156 22484 16212 23102
rect 16828 23042 16884 23324
rect 16828 22990 16830 23042
rect 16882 22990 16884 23042
rect 16268 22932 16324 22942
rect 16268 22838 16324 22876
rect 15932 22370 15988 22428
rect 15932 22318 15934 22370
rect 15986 22318 15988 22370
rect 15932 22306 15988 22318
rect 16044 22482 16212 22484
rect 16044 22430 16158 22482
rect 16210 22430 16212 22482
rect 16044 22428 16212 22430
rect 16044 22036 16100 22428
rect 16156 22418 16212 22428
rect 16604 22260 16660 22270
rect 16604 22166 16660 22204
rect 15820 21980 16100 22036
rect 15820 21700 15876 21980
rect 15260 21698 15876 21700
rect 15260 21646 15822 21698
rect 15874 21646 15876 21698
rect 15260 21644 15876 21646
rect 15260 21586 15316 21644
rect 15820 21634 15876 21644
rect 16492 21700 16548 21710
rect 15260 21534 15262 21586
rect 15314 21534 15316 21586
rect 15260 21522 15316 21534
rect 15932 21586 15988 21598
rect 15932 21534 15934 21586
rect 15986 21534 15988 21586
rect 15484 21476 15540 21486
rect 15372 21474 15540 21476
rect 15372 21422 15486 21474
rect 15538 21422 15540 21474
rect 15372 21420 15540 21422
rect 15372 20802 15428 21420
rect 15484 21410 15540 21420
rect 15932 21028 15988 21534
rect 16492 21586 16548 21644
rect 16828 21700 16884 22990
rect 16828 21634 16884 21644
rect 16492 21534 16494 21586
rect 16546 21534 16548 21586
rect 16492 21522 16548 21534
rect 15932 20962 15988 20972
rect 15372 20750 15374 20802
rect 15426 20750 15428 20802
rect 15372 19908 15428 20750
rect 15708 20916 15764 20926
rect 15708 20802 15764 20860
rect 16492 20804 16548 20814
rect 15708 20750 15710 20802
rect 15762 20750 15764 20802
rect 15708 20738 15764 20750
rect 16380 20802 16548 20804
rect 16380 20750 16494 20802
rect 16546 20750 16548 20802
rect 16380 20748 16548 20750
rect 15820 20690 15876 20702
rect 15820 20638 15822 20690
rect 15874 20638 15876 20690
rect 15820 20132 15876 20638
rect 15820 20066 15876 20076
rect 16044 20580 16100 20590
rect 15372 19852 15988 19908
rect 15148 19628 15316 19684
rect 15260 19572 15316 19628
rect 15260 19516 15540 19572
rect 15148 19460 15204 19470
rect 15036 19348 15092 19358
rect 15036 18674 15092 19292
rect 15148 19346 15204 19404
rect 15148 19294 15150 19346
rect 15202 19294 15204 19346
rect 15148 19282 15204 19294
rect 15372 19348 15428 19358
rect 15036 18622 15038 18674
rect 15090 18622 15092 18674
rect 15036 18610 15092 18622
rect 15260 19234 15316 19246
rect 15260 19182 15262 19234
rect 15314 19182 15316 19234
rect 14924 18510 14926 18562
rect 14978 18510 14980 18562
rect 14924 18498 14980 18510
rect 15260 18452 15316 19182
rect 15260 18358 15316 18396
rect 15372 18450 15428 19292
rect 15372 18398 15374 18450
rect 15426 18398 15428 18450
rect 15372 18386 15428 18398
rect 14364 18228 14420 18238
rect 14252 17892 14308 17902
rect 14140 17780 14196 17790
rect 14140 17686 14196 17724
rect 14252 17778 14308 17836
rect 14252 17726 14254 17778
rect 14306 17726 14308 17778
rect 14252 17714 14308 17726
rect 14364 17556 14420 18172
rect 14364 17462 14420 17500
rect 14700 17780 14756 17790
rect 14028 17378 14084 17388
rect 14140 17108 14196 17118
rect 13244 17042 13300 17052
rect 13804 17106 14196 17108
rect 13804 17054 14142 17106
rect 14194 17054 14196 17106
rect 13804 17052 14196 17054
rect 13804 16996 13860 17052
rect 12796 16830 12798 16882
rect 12850 16830 12852 16882
rect 12796 16322 12852 16830
rect 13356 16940 13860 16996
rect 13356 16882 13412 16940
rect 13356 16830 13358 16882
rect 13410 16830 13412 16882
rect 13356 16818 13412 16830
rect 12796 16270 12798 16322
rect 12850 16270 12852 16322
rect 12796 16258 12852 16270
rect 13468 16324 13524 16334
rect 13468 16230 13524 16268
rect 13580 16212 13636 16940
rect 13916 16884 13972 16894
rect 13916 16790 13972 16828
rect 13580 16118 13636 16156
rect 12572 15934 12574 15986
rect 12626 15934 12628 15986
rect 12572 15922 12628 15934
rect 13580 15540 13636 15550
rect 13580 15446 13636 15484
rect 14140 15538 14196 17052
rect 14252 16996 14308 17006
rect 14252 16902 14308 16940
rect 14140 15486 14142 15538
rect 14194 15486 14196 15538
rect 14140 15474 14196 15486
rect 14252 16212 14308 16222
rect 14700 16212 14756 17724
rect 15372 17668 15428 17678
rect 14924 17556 14980 17566
rect 14924 17462 14980 17500
rect 15372 17444 15428 17612
rect 15372 17350 15428 17388
rect 15484 17106 15540 19516
rect 15820 19460 15876 19470
rect 15820 18562 15876 19404
rect 15932 19346 15988 19852
rect 15932 19294 15934 19346
rect 15986 19294 15988 19346
rect 15932 19282 15988 19294
rect 16044 19348 16100 20524
rect 16044 19282 16100 19292
rect 16380 20468 16436 20748
rect 16492 20738 16548 20748
rect 15932 18676 15988 18686
rect 16380 18676 16436 20412
rect 16716 20130 16772 20142
rect 16716 20078 16718 20130
rect 16770 20078 16772 20130
rect 16716 20020 16772 20078
rect 16716 19954 16772 19964
rect 16940 19796 16996 26908
rect 17164 25956 17220 28364
rect 17724 28082 17780 28812
rect 17836 28866 17892 29596
rect 17948 29652 18004 29662
rect 18060 29652 18116 30828
rect 18172 30322 18228 30940
rect 18620 30884 18676 31726
rect 18732 31556 18788 31566
rect 18732 31462 18788 31500
rect 18844 31554 18900 33068
rect 18844 31502 18846 31554
rect 18898 31502 18900 31554
rect 18172 30270 18174 30322
rect 18226 30270 18228 30322
rect 18172 30258 18228 30270
rect 18284 30828 18676 30884
rect 18732 30994 18788 31006
rect 18732 30942 18734 30994
rect 18786 30942 18788 30994
rect 18732 30884 18788 30942
rect 18284 30434 18340 30828
rect 18732 30818 18788 30828
rect 18844 30660 18900 31502
rect 18956 31220 19012 34300
rect 19180 34244 19236 34254
rect 19292 34244 19348 35084
rect 19404 35026 19460 35644
rect 19404 34974 19406 35026
rect 19458 34974 19460 35026
rect 19404 34962 19460 34974
rect 19516 34244 19572 35756
rect 19628 35718 19684 35756
rect 19740 35700 19796 35710
rect 20188 35700 20244 36206
rect 20412 36260 20468 36270
rect 20412 36166 20468 36204
rect 20972 36260 21028 36270
rect 20412 36036 20468 36046
rect 19796 35644 20244 35700
rect 20300 35700 20356 35710
rect 19740 35606 19796 35644
rect 20300 35586 20356 35644
rect 20300 35534 20302 35586
rect 20354 35534 20356 35586
rect 19852 35364 19908 35374
rect 19852 35026 19908 35308
rect 19852 34974 19854 35026
rect 19906 34974 19908 35026
rect 19852 34962 19908 34974
rect 20300 34804 20356 35534
rect 20412 35026 20468 35980
rect 20748 35588 20804 35598
rect 20748 35494 20804 35532
rect 20972 35364 21028 36204
rect 21308 36258 21364 36270
rect 21308 36206 21310 36258
rect 21362 36206 21364 36258
rect 21308 35924 21364 36206
rect 21532 36260 21588 36298
rect 21532 36194 21588 36204
rect 21532 36036 21588 36046
rect 21644 36036 21700 38612
rect 22092 38052 22148 38062
rect 21868 38050 22148 38052
rect 21868 37998 22094 38050
rect 22146 37998 22148 38050
rect 21868 37996 22148 37998
rect 21588 35980 21700 36036
rect 21756 36372 21812 36382
rect 21532 35970 21588 35980
rect 21420 35924 21476 35934
rect 21756 35924 21812 36316
rect 21308 35922 21476 35924
rect 21308 35870 21422 35922
rect 21474 35870 21476 35922
rect 21308 35868 21476 35870
rect 21420 35858 21476 35868
rect 21644 35868 21812 35924
rect 20972 35298 21028 35308
rect 21084 35698 21140 35710
rect 21084 35646 21086 35698
rect 21138 35646 21140 35698
rect 20748 35140 20804 35150
rect 20748 35046 20804 35084
rect 20412 34974 20414 35026
rect 20466 34974 20468 35026
rect 20412 34962 20468 34974
rect 20636 35028 20692 35038
rect 20300 34738 20356 34748
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19292 34188 19460 34244
rect 19516 34188 19684 34244
rect 19180 34130 19236 34188
rect 19180 34078 19182 34130
rect 19234 34078 19236 34130
rect 19180 34066 19236 34078
rect 19404 34020 19460 34188
rect 19516 34020 19572 34030
rect 19404 34018 19572 34020
rect 19404 33966 19518 34018
rect 19570 33966 19572 34018
rect 19404 33964 19572 33966
rect 19068 33460 19124 33470
rect 19068 33366 19124 33404
rect 19180 33124 19236 33134
rect 19180 33030 19236 33068
rect 19404 33124 19460 33134
rect 19404 33030 19460 33068
rect 19292 32676 19348 32686
rect 19292 32582 19348 32620
rect 19404 32564 19460 32574
rect 19404 32470 19460 32508
rect 19404 31892 19460 31902
rect 19180 31890 19460 31892
rect 19180 31838 19406 31890
rect 19458 31838 19460 31890
rect 19180 31836 19460 31838
rect 18956 31164 19124 31220
rect 18956 30996 19012 31006
rect 18956 30902 19012 30940
rect 18284 30382 18286 30434
rect 18338 30382 18340 30434
rect 18284 30212 18340 30382
rect 18508 30604 18900 30660
rect 18508 30324 18564 30604
rect 19068 30548 19124 31164
rect 18844 30492 19124 30548
rect 19180 30882 19236 31836
rect 19404 31826 19460 31836
rect 19516 31780 19572 33964
rect 19628 32004 19684 34188
rect 20636 34130 20692 34972
rect 20636 34078 20638 34130
rect 20690 34078 20692 34130
rect 20636 34066 20692 34078
rect 20972 34916 21028 34926
rect 20972 34130 21028 34860
rect 21084 34242 21140 35646
rect 21308 35700 21364 35710
rect 21308 35364 21364 35644
rect 21308 35298 21364 35308
rect 21532 35698 21588 35710
rect 21532 35646 21534 35698
rect 21586 35646 21588 35698
rect 21084 34190 21086 34242
rect 21138 34190 21140 34242
rect 21084 34178 21140 34190
rect 21420 34244 21476 34254
rect 21532 34244 21588 35646
rect 21420 34242 21588 34244
rect 21420 34190 21422 34242
rect 21474 34190 21588 34242
rect 21420 34188 21588 34190
rect 21420 34178 21476 34188
rect 20972 34078 20974 34130
rect 21026 34078 21028 34130
rect 19964 33124 20020 33162
rect 19964 33058 20020 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20188 32452 20244 32462
rect 19628 31948 19796 32004
rect 19516 31714 19572 31724
rect 19180 30830 19182 30882
rect 19234 30830 19236 30882
rect 18508 30258 18564 30268
rect 18620 30436 18676 30446
rect 18284 30146 18340 30156
rect 18620 30210 18676 30380
rect 18620 30158 18622 30210
rect 18674 30158 18676 30210
rect 18004 29596 18116 29652
rect 18172 30100 18228 30110
rect 17948 29586 18004 29596
rect 18172 29426 18228 30044
rect 18172 29374 18174 29426
rect 18226 29374 18228 29426
rect 18172 29362 18228 29374
rect 18620 29426 18676 30158
rect 18620 29374 18622 29426
rect 18674 29374 18676 29426
rect 18620 29362 18676 29374
rect 18732 30212 18788 30222
rect 17836 28814 17838 28866
rect 17890 28814 17892 28866
rect 17836 28802 17892 28814
rect 17948 28756 18004 28766
rect 17948 28662 18004 28700
rect 18620 28756 18676 28766
rect 18396 28420 18452 28430
rect 18396 28326 18452 28364
rect 17724 28030 17726 28082
rect 17778 28030 17780 28082
rect 17388 26964 17444 27002
rect 17388 26898 17444 26908
rect 17724 26516 17780 28030
rect 18284 28084 18340 28094
rect 18284 27412 18340 28028
rect 18284 27356 18564 27412
rect 18284 27074 18340 27356
rect 18284 27022 18286 27074
rect 18338 27022 18340 27074
rect 18284 27010 18340 27022
rect 18396 27188 18452 27198
rect 18396 26908 18452 27132
rect 17724 26450 17780 26460
rect 17948 26852 18004 26862
rect 17948 26178 18004 26796
rect 17948 26126 17950 26178
rect 18002 26126 18004 26178
rect 17948 26114 18004 26126
rect 18284 26852 18452 26908
rect 17164 25900 17668 25956
rect 17052 25508 17108 25518
rect 17052 22370 17108 25452
rect 17276 25506 17332 25518
rect 17276 25454 17278 25506
rect 17330 25454 17332 25506
rect 17276 24948 17332 25454
rect 17276 24882 17332 24892
rect 17500 24834 17556 24846
rect 17500 24782 17502 24834
rect 17554 24782 17556 24834
rect 17388 24724 17444 24734
rect 17388 24630 17444 24668
rect 17500 24612 17556 24782
rect 17500 24546 17556 24556
rect 17612 24388 17668 25900
rect 18060 25060 18116 25070
rect 17500 24332 17668 24388
rect 17724 24722 17780 24734
rect 17724 24670 17726 24722
rect 17778 24670 17780 24722
rect 17276 23604 17332 23614
rect 17164 23492 17332 23548
rect 17500 23492 17556 24332
rect 17724 23548 17780 24670
rect 18060 24610 18116 25004
rect 18060 24558 18062 24610
rect 18114 24558 18116 24610
rect 17948 24498 18004 24510
rect 17948 24446 17950 24498
rect 18002 24446 18004 24498
rect 17836 23716 17892 23726
rect 17948 23716 18004 24446
rect 18060 23828 18116 24558
rect 18060 23762 18116 23772
rect 17836 23714 18004 23716
rect 17836 23662 17838 23714
rect 17890 23662 18004 23714
rect 17836 23660 18004 23662
rect 17836 23650 17892 23660
rect 17724 23492 17892 23548
rect 17164 23156 17220 23492
rect 17500 23436 17668 23492
rect 17836 23436 18004 23492
rect 17612 23380 17668 23436
rect 17612 23324 17892 23380
rect 17500 23268 17556 23278
rect 17500 23174 17556 23212
rect 17612 23212 17780 23268
rect 17164 23100 17332 23156
rect 17052 22318 17054 22370
rect 17106 22318 17108 22370
rect 17052 21476 17108 22318
rect 17164 22260 17220 22270
rect 17164 22166 17220 22204
rect 17052 21410 17108 21420
rect 17052 20804 17108 20814
rect 17276 20804 17332 23100
rect 17388 23154 17444 23166
rect 17388 23102 17390 23154
rect 17442 23102 17444 23154
rect 17388 22482 17444 23102
rect 17612 23154 17668 23212
rect 17612 23102 17614 23154
rect 17666 23102 17668 23154
rect 17612 23090 17668 23102
rect 17724 23156 17780 23212
rect 17724 23090 17780 23100
rect 17388 22430 17390 22482
rect 17442 22430 17444 22482
rect 17388 22418 17444 22430
rect 17612 22370 17668 22382
rect 17612 22318 17614 22370
rect 17666 22318 17668 22370
rect 17388 22148 17444 22158
rect 17388 22054 17444 22092
rect 17500 21812 17556 21822
rect 17500 21718 17556 21756
rect 17612 21810 17668 22318
rect 17612 21758 17614 21810
rect 17666 21758 17668 21810
rect 17612 21746 17668 21758
rect 17724 21812 17780 21822
rect 17836 21812 17892 23324
rect 17948 23154 18004 23436
rect 17948 23102 17950 23154
rect 18002 23102 18004 23154
rect 17948 23090 18004 23102
rect 18060 22932 18116 22942
rect 18060 22370 18116 22876
rect 18060 22318 18062 22370
rect 18114 22318 18116 22370
rect 18060 22306 18116 22318
rect 18172 22148 18228 22158
rect 18172 22054 18228 22092
rect 17780 21756 17892 21812
rect 17948 22036 18004 22046
rect 17724 21746 17780 21756
rect 17948 21700 18004 21980
rect 18284 21700 18340 26852
rect 18508 26290 18564 27356
rect 18620 26908 18676 28700
rect 18732 27188 18788 30156
rect 18732 27122 18788 27132
rect 18620 26852 18788 26908
rect 18508 26238 18510 26290
rect 18562 26238 18564 26290
rect 18508 26180 18564 26238
rect 18620 26180 18676 26190
rect 18508 26178 18676 26180
rect 18508 26126 18622 26178
rect 18674 26126 18676 26178
rect 18508 26124 18676 26126
rect 18508 23828 18564 26124
rect 18620 26114 18676 26124
rect 18732 25172 18788 26852
rect 18844 25732 18900 30492
rect 19180 30436 19236 30830
rect 19180 30370 19236 30380
rect 19292 31668 19348 31678
rect 19292 30324 19348 31612
rect 19740 31668 19796 31948
rect 19740 31602 19796 31612
rect 19516 31556 19572 31566
rect 19572 31500 19684 31556
rect 19516 31490 19572 31500
rect 19516 31220 19572 31230
rect 19516 31126 19572 31164
rect 19628 31108 19684 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20188 31220 20244 32396
rect 20972 32452 21028 34078
rect 20972 32358 21028 32396
rect 20076 31164 20244 31220
rect 20524 31780 20580 31790
rect 19628 31052 20020 31108
rect 19404 30996 19460 31006
rect 19404 30994 19572 30996
rect 19404 30942 19406 30994
rect 19458 30942 19572 30994
rect 19404 30940 19572 30942
rect 19404 30930 19460 30940
rect 19404 30324 19460 30334
rect 19292 30322 19460 30324
rect 19292 30270 19406 30322
rect 19458 30270 19460 30322
rect 19292 30268 19460 30270
rect 19404 30258 19460 30268
rect 19180 30210 19236 30222
rect 19180 30158 19182 30210
rect 19234 30158 19236 30210
rect 19180 29652 19236 30158
rect 19404 29988 19460 29998
rect 19292 29652 19348 29662
rect 19180 29596 19292 29652
rect 19292 29586 19348 29596
rect 19404 29650 19460 29932
rect 19516 29764 19572 30940
rect 19964 30994 20020 31052
rect 19964 30942 19966 30994
rect 20018 30942 20020 30994
rect 19964 30930 20020 30942
rect 19740 30882 19796 30894
rect 19740 30830 19742 30882
rect 19794 30830 19796 30882
rect 19740 30772 19796 30830
rect 20076 30772 20132 31164
rect 20524 30884 20580 31724
rect 20748 31780 20804 31790
rect 20636 31220 20692 31230
rect 20636 31106 20692 31164
rect 20748 31218 20804 31724
rect 20748 31166 20750 31218
rect 20802 31166 20804 31218
rect 20748 31154 20804 31166
rect 20636 31054 20638 31106
rect 20690 31054 20692 31106
rect 20636 31042 20692 31054
rect 20972 30996 21028 31006
rect 20972 30994 21476 30996
rect 20972 30942 20974 30994
rect 21026 30942 21476 30994
rect 20972 30940 21476 30942
rect 20972 30930 21028 30940
rect 20524 30828 20692 30884
rect 19740 30716 20132 30772
rect 20300 30772 20356 30782
rect 20300 30770 20580 30772
rect 20300 30718 20302 30770
rect 20354 30718 20580 30770
rect 20300 30716 20580 30718
rect 20300 30706 20356 30716
rect 20076 30212 20132 30222
rect 20076 30118 20132 30156
rect 20524 30210 20580 30716
rect 20524 30158 20526 30210
rect 20578 30158 20580 30210
rect 20524 30146 20580 30158
rect 20412 30098 20468 30110
rect 20412 30046 20414 30098
rect 20466 30046 20468 30098
rect 20188 29986 20244 29998
rect 20188 29934 20190 29986
rect 20242 29934 20244 29986
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19516 29698 19572 29708
rect 19404 29598 19406 29650
rect 19458 29598 19460 29650
rect 19404 29586 19460 29598
rect 19068 29540 19124 29550
rect 19068 29446 19124 29484
rect 20188 29540 20244 29934
rect 20300 29988 20356 29998
rect 20412 29988 20468 30046
rect 20524 29988 20580 29998
rect 20412 29932 20524 29988
rect 20300 29894 20356 29932
rect 20524 29922 20580 29932
rect 20412 29652 20468 29662
rect 20412 29558 20468 29596
rect 20188 29474 20244 29484
rect 19516 29426 19572 29438
rect 19516 29374 19518 29426
rect 19570 29374 19572 29426
rect 19068 28420 19124 28430
rect 19180 28420 19236 28430
rect 19068 28418 19180 28420
rect 19068 28366 19070 28418
rect 19122 28366 19180 28418
rect 19068 28364 19180 28366
rect 19068 28354 19124 28364
rect 19068 27860 19124 27870
rect 19068 27766 19124 27804
rect 19068 27076 19124 27086
rect 18956 26852 19012 26862
rect 19068 26852 19124 27020
rect 18956 26850 19124 26852
rect 18956 26798 18958 26850
rect 19010 26798 19124 26850
rect 18956 26796 19124 26798
rect 19180 26852 19236 28364
rect 19516 27858 19572 29374
rect 19628 29426 19684 29438
rect 19628 29374 19630 29426
rect 19682 29374 19684 29426
rect 19628 28420 19684 29374
rect 19964 29428 20020 29438
rect 19964 28756 20020 29372
rect 20076 29426 20132 29438
rect 20076 29374 20078 29426
rect 20130 29374 20132 29426
rect 20076 29204 20132 29374
rect 20300 29428 20356 29438
rect 20636 29428 20692 30828
rect 21308 30436 21364 30446
rect 21308 30342 21364 30380
rect 21420 30322 21476 30940
rect 21644 30436 21700 35868
rect 21756 35700 21812 35710
rect 21756 35606 21812 35644
rect 21868 35252 21924 37996
rect 22092 37986 22148 37996
rect 22204 37604 22260 41200
rect 22876 38162 22932 41200
rect 23548 38668 23604 41200
rect 24220 39620 24276 41200
rect 24220 39564 24836 39620
rect 23548 38612 23716 38668
rect 22876 38110 22878 38162
rect 22930 38110 22932 38162
rect 22876 38098 22932 38110
rect 23436 38052 23492 38062
rect 22204 37538 22260 37548
rect 23212 38050 23492 38052
rect 23212 37998 23438 38050
rect 23490 37998 23492 38050
rect 23212 37996 23492 37998
rect 22652 37492 22708 37502
rect 23212 37492 23268 37996
rect 23436 37986 23492 37996
rect 22652 37490 22932 37492
rect 22652 37438 22654 37490
rect 22706 37438 22932 37490
rect 22652 37436 22932 37438
rect 22652 37426 22708 37436
rect 22876 36706 22932 37436
rect 22876 36654 22878 36706
rect 22930 36654 22932 36706
rect 22876 36642 22932 36654
rect 23100 37490 23268 37492
rect 23100 37438 23214 37490
rect 23266 37438 23268 37490
rect 23100 37436 23268 37438
rect 21980 36482 22036 36494
rect 21980 36430 21982 36482
rect 22034 36430 22036 36482
rect 21980 35922 22036 36430
rect 22316 36428 22708 36484
rect 22204 36260 22260 36270
rect 22092 36258 22260 36260
rect 22092 36206 22206 36258
rect 22258 36206 22260 36258
rect 22092 36204 22260 36206
rect 22092 36036 22148 36204
rect 22204 36194 22260 36204
rect 22092 35970 22148 35980
rect 21980 35870 21982 35922
rect 22034 35870 22036 35922
rect 21980 35858 22036 35870
rect 22204 35924 22260 35934
rect 22316 35924 22372 36428
rect 22204 35922 22372 35924
rect 22204 35870 22206 35922
rect 22258 35870 22372 35922
rect 22204 35868 22372 35870
rect 22540 36258 22596 36270
rect 22540 36206 22542 36258
rect 22594 36206 22596 36258
rect 21868 35196 22148 35252
rect 21980 35028 22036 35038
rect 21756 34916 21812 34926
rect 21756 33346 21812 34860
rect 21756 33294 21758 33346
rect 21810 33294 21812 33346
rect 21756 33282 21812 33294
rect 21980 33346 22036 34972
rect 22092 34356 22148 35196
rect 22204 34914 22260 35868
rect 22316 35698 22372 35710
rect 22316 35646 22318 35698
rect 22370 35646 22372 35698
rect 22316 35588 22372 35646
rect 22316 35522 22372 35532
rect 22204 34862 22206 34914
rect 22258 34862 22260 34914
rect 22204 34850 22260 34862
rect 22428 35028 22484 35038
rect 22428 34914 22484 34972
rect 22428 34862 22430 34914
rect 22482 34862 22484 34914
rect 22428 34850 22484 34862
rect 22428 34468 22484 34478
rect 22092 34300 22260 34356
rect 21980 33294 21982 33346
rect 22034 33294 22036 33346
rect 21980 33282 22036 33294
rect 22092 34130 22148 34142
rect 22092 34078 22094 34130
rect 22146 34078 22148 34130
rect 22092 34020 22148 34078
rect 21868 33236 21924 33274
rect 21868 33170 21924 33180
rect 21980 33124 22036 33134
rect 21420 30270 21422 30322
rect 21474 30270 21476 30322
rect 21420 30258 21476 30270
rect 21532 30380 21700 30436
rect 21868 32452 21924 32462
rect 20356 29372 20692 29428
rect 20972 29988 21028 29998
rect 20300 29334 20356 29372
rect 20972 29316 21028 29932
rect 20972 29222 21028 29260
rect 20412 29204 20468 29214
rect 20076 29202 20468 29204
rect 20076 29150 20414 29202
rect 20466 29150 20468 29202
rect 20076 29148 20468 29150
rect 20412 29138 20468 29148
rect 19964 28662 20020 28700
rect 21420 28756 21476 28766
rect 21532 28756 21588 30380
rect 21644 30212 21700 30222
rect 21868 30212 21924 32396
rect 21980 32004 22036 33068
rect 22092 32228 22148 33964
rect 22204 32452 22260 34300
rect 22316 34132 22372 34142
rect 22316 34038 22372 34076
rect 22428 33346 22484 34412
rect 22428 33294 22430 33346
rect 22482 33294 22484 33346
rect 22428 33282 22484 33294
rect 22204 32386 22260 32396
rect 22428 32228 22484 32238
rect 22092 32172 22428 32228
rect 22428 32162 22484 32172
rect 21980 31938 22036 31948
rect 22204 31778 22260 31790
rect 22204 31726 22206 31778
rect 22258 31726 22260 31778
rect 22204 31668 22260 31726
rect 22428 31780 22484 31790
rect 22428 31686 22484 31724
rect 21644 30210 21924 30212
rect 21644 30158 21646 30210
rect 21698 30158 21924 30210
rect 21644 30156 21924 30158
rect 22092 30212 22148 30222
rect 21644 29652 21700 30156
rect 22092 29986 22148 30156
rect 22204 30100 22260 31612
rect 22540 31220 22596 36206
rect 22652 36148 22708 36428
rect 22988 36372 23044 36382
rect 22988 36278 23044 36316
rect 23100 36148 23156 37436
rect 23212 37426 23268 37436
rect 23548 37268 23604 37278
rect 22652 36092 23156 36148
rect 23436 37154 23492 37166
rect 23436 37102 23438 37154
rect 23490 37102 23492 37154
rect 22764 35922 22820 36092
rect 22764 35870 22766 35922
rect 22818 35870 22820 35922
rect 22764 35858 22820 35870
rect 22652 35698 22708 35710
rect 22652 35646 22654 35698
rect 22706 35646 22708 35698
rect 22652 35140 22708 35646
rect 22652 35074 22708 35084
rect 22764 35474 22820 35486
rect 22764 35422 22766 35474
rect 22818 35422 22820 35474
rect 22652 34802 22708 34814
rect 22652 34750 22654 34802
rect 22706 34750 22708 34802
rect 22652 34132 22708 34750
rect 22764 34244 22820 35422
rect 23436 35140 23492 37102
rect 23548 36482 23604 37212
rect 23660 36820 23716 38612
rect 24780 38162 24836 39564
rect 25564 38610 25620 41200
rect 25564 38558 25566 38610
rect 25618 38558 25620 38610
rect 25564 38546 25620 38558
rect 26236 38612 26292 41200
rect 26908 38836 26964 41200
rect 26908 38780 27188 38836
rect 26236 38546 26292 38556
rect 26348 38610 26404 38622
rect 27020 38612 27076 38622
rect 26348 38558 26350 38610
rect 26402 38558 26404 38610
rect 24780 38110 24782 38162
rect 24834 38110 24836 38162
rect 24780 38098 24836 38110
rect 26348 38162 26404 38558
rect 26348 38110 26350 38162
rect 26402 38110 26404 38162
rect 26348 38098 26404 38110
rect 26908 38610 27076 38612
rect 26908 38558 27022 38610
rect 27074 38558 27076 38610
rect 26908 38556 27076 38558
rect 25564 38052 25620 38062
rect 25452 38050 25620 38052
rect 25452 37998 25566 38050
rect 25618 37998 25620 38050
rect 25452 37996 25620 37998
rect 23996 37828 24052 37838
rect 23660 36754 23716 36764
rect 23884 37826 24052 37828
rect 23884 37774 23998 37826
rect 24050 37774 24052 37826
rect 23884 37772 24052 37774
rect 23548 36430 23550 36482
rect 23602 36430 23604 36482
rect 23548 36418 23604 36430
rect 23884 36372 23940 37772
rect 23996 37762 24052 37772
rect 23996 37604 24052 37614
rect 23996 37490 24052 37548
rect 23996 37438 23998 37490
rect 24050 37438 24052 37490
rect 23996 37426 24052 37438
rect 24332 37380 24388 37390
rect 23884 36306 23940 36316
rect 24108 37378 24388 37380
rect 24108 37326 24334 37378
rect 24386 37326 24388 37378
rect 24108 37324 24388 37326
rect 24108 36036 24164 37324
rect 24332 37314 24388 37324
rect 25228 37380 25284 37390
rect 25228 37286 25284 37324
rect 25340 37378 25396 37390
rect 25340 37326 25342 37378
rect 25394 37326 25396 37378
rect 24668 37266 24724 37278
rect 24668 37214 24670 37266
rect 24722 37214 24724 37266
rect 24668 36820 24724 37214
rect 25340 37044 25396 37326
rect 24668 36754 24724 36764
rect 25116 36988 25340 37044
rect 24220 36484 24276 36494
rect 24220 36390 24276 36428
rect 22988 35084 23492 35140
rect 23548 35980 24164 36036
rect 23548 35810 23604 35980
rect 23548 35758 23550 35810
rect 23602 35758 23604 35810
rect 22988 35028 23044 35084
rect 22988 34934 23044 34972
rect 23212 34914 23268 34926
rect 23212 34862 23214 34914
rect 23266 34862 23268 34914
rect 23212 34692 23268 34862
rect 23436 34916 23492 34926
rect 23436 34822 23492 34860
rect 23548 34692 23604 35758
rect 23212 34636 23604 34692
rect 23660 35810 23716 35822
rect 23660 35758 23662 35810
rect 23714 35758 23716 35810
rect 23436 34468 23492 34636
rect 22764 34178 22820 34188
rect 23324 34356 23380 34366
rect 22652 32674 22708 34076
rect 23324 34130 23380 34300
rect 23324 34078 23326 34130
rect 23378 34078 23380 34130
rect 23324 34066 23380 34078
rect 23436 34018 23492 34412
rect 23660 34356 23716 35758
rect 24668 35812 24724 35822
rect 25116 35812 25172 36988
rect 25340 36950 25396 36988
rect 25340 36484 25396 36494
rect 25340 35922 25396 36428
rect 25340 35870 25342 35922
rect 25394 35870 25396 35922
rect 25340 35858 25396 35870
rect 25452 35924 25508 37996
rect 25564 37986 25620 37996
rect 25788 37380 25844 37390
rect 25564 37268 25620 37278
rect 25564 37266 25732 37268
rect 25564 37214 25566 37266
rect 25618 37214 25732 37266
rect 25564 37212 25732 37214
rect 25564 37202 25620 37212
rect 25452 35868 25620 35924
rect 24668 35810 25172 35812
rect 24668 35758 24670 35810
rect 24722 35758 25172 35810
rect 24668 35756 25172 35758
rect 24668 35746 24724 35756
rect 23884 35700 23940 35710
rect 24220 35700 24276 35710
rect 23884 35698 24052 35700
rect 23884 35646 23886 35698
rect 23938 35646 24052 35698
rect 23884 35644 24052 35646
rect 23884 35634 23940 35644
rect 23996 35474 24052 35644
rect 23996 35422 23998 35474
rect 24050 35422 24052 35474
rect 23996 35410 24052 35422
rect 24220 34916 24276 35644
rect 25228 35698 25284 35710
rect 25228 35646 25230 35698
rect 25282 35646 25284 35698
rect 24332 35476 24388 35486
rect 24332 35474 24500 35476
rect 24332 35422 24334 35474
rect 24386 35422 24500 35474
rect 24332 35420 24500 35422
rect 24332 35410 24388 35420
rect 24332 35252 24388 35262
rect 24444 35252 24500 35420
rect 24556 35474 24612 35486
rect 24556 35422 24558 35474
rect 24610 35422 24612 35474
rect 24556 35364 24612 35422
rect 24556 35308 25172 35364
rect 24444 35196 25060 35252
rect 24332 34916 24388 35196
rect 24556 35028 24612 35038
rect 24556 34934 24612 34972
rect 24332 34860 24500 34916
rect 24220 34822 24276 34860
rect 24444 34804 24500 34860
rect 24556 34804 24612 34814
rect 24444 34748 24556 34804
rect 24556 34710 24612 34748
rect 23660 34290 23716 34300
rect 23884 34690 23940 34702
rect 23884 34638 23886 34690
rect 23938 34638 23940 34690
rect 23772 34020 23828 34030
rect 23436 33966 23438 34018
rect 23490 33966 23492 34018
rect 23436 33954 23492 33966
rect 23548 34018 23828 34020
rect 23548 33966 23774 34018
rect 23826 33966 23828 34018
rect 23548 33964 23828 33966
rect 23548 33796 23604 33964
rect 23772 33954 23828 33964
rect 23884 33908 23940 34638
rect 24332 34692 24388 34702
rect 24332 34690 24500 34692
rect 24332 34638 24334 34690
rect 24386 34638 24500 34690
rect 24332 34636 24500 34638
rect 24332 34626 24388 34636
rect 24108 34132 24164 34142
rect 24108 34038 24164 34076
rect 24332 34130 24388 34142
rect 24332 34078 24334 34130
rect 24386 34078 24388 34130
rect 24220 34018 24276 34030
rect 24220 33966 24222 34018
rect 24274 33966 24276 34018
rect 23996 33908 24052 33918
rect 23884 33852 23996 33908
rect 23996 33842 24052 33852
rect 23436 33740 23604 33796
rect 23436 33460 23492 33740
rect 24220 33684 24276 33966
rect 24332 34020 24388 34078
rect 24332 33954 24388 33964
rect 23212 33404 23492 33460
rect 23548 33628 24276 33684
rect 23212 33346 23268 33404
rect 23212 33294 23214 33346
rect 23266 33294 23268 33346
rect 23212 33282 23268 33294
rect 23324 32786 23380 33404
rect 23548 33346 23604 33628
rect 24444 33572 24500 34636
rect 24668 34690 24724 34702
rect 24668 34638 24670 34690
rect 24722 34638 24724 34690
rect 24668 34356 24724 34638
rect 24780 34468 24836 34478
rect 24836 34412 24948 34468
rect 24780 34402 24836 34412
rect 23660 33516 24500 33572
rect 24556 34300 24724 34356
rect 24556 33570 24612 34300
rect 24668 34132 24724 34142
rect 24668 34038 24724 34076
rect 24892 34132 24948 34412
rect 24892 34066 24948 34076
rect 24556 33518 24558 33570
rect 24610 33518 24612 33570
rect 23660 33458 23716 33516
rect 24556 33506 24612 33518
rect 23660 33406 23662 33458
rect 23714 33406 23716 33458
rect 23660 33394 23716 33406
rect 23548 33294 23550 33346
rect 23602 33294 23604 33346
rect 23548 33282 23604 33294
rect 23996 33348 24052 33358
rect 23996 33254 24052 33292
rect 24220 33346 24276 33358
rect 24220 33294 24222 33346
rect 24274 33294 24276 33346
rect 24220 33236 24276 33294
rect 24220 33170 24276 33180
rect 25004 33234 25060 35196
rect 25116 34356 25172 35308
rect 25228 35028 25284 35646
rect 25452 35698 25508 35710
rect 25452 35646 25454 35698
rect 25506 35646 25508 35698
rect 25452 35138 25508 35646
rect 25452 35086 25454 35138
rect 25506 35086 25508 35138
rect 25452 35074 25508 35086
rect 25228 34962 25284 34972
rect 25228 34804 25284 34814
rect 25228 34710 25284 34748
rect 25452 34356 25508 34366
rect 25172 34354 25508 34356
rect 25172 34302 25454 34354
rect 25506 34302 25508 34354
rect 25172 34300 25508 34302
rect 25116 34262 25172 34300
rect 25452 34290 25508 34300
rect 25228 34132 25284 34142
rect 25228 34038 25284 34076
rect 25340 34018 25396 34030
rect 25340 33966 25342 34018
rect 25394 33966 25396 34018
rect 25340 33572 25396 33966
rect 25116 33516 25396 33572
rect 25116 33346 25172 33516
rect 25116 33294 25118 33346
rect 25170 33294 25172 33346
rect 25116 33282 25172 33294
rect 25004 33182 25006 33234
rect 25058 33182 25060 33234
rect 25004 33170 25060 33182
rect 23324 32734 23326 32786
rect 23378 32734 23380 32786
rect 23324 32722 23380 32734
rect 24780 33122 24836 33134
rect 24780 33070 24782 33122
rect 24834 33070 24836 33122
rect 22652 32622 22654 32674
rect 22706 32622 22708 32674
rect 22652 32610 22708 32622
rect 24108 32676 24164 32686
rect 24108 32582 24164 32620
rect 22764 32564 22820 32574
rect 23212 32564 23268 32574
rect 22764 32562 23268 32564
rect 22764 32510 22766 32562
rect 22818 32510 23214 32562
rect 23266 32510 23268 32562
rect 22764 32508 23268 32510
rect 22764 32498 22820 32508
rect 23212 32498 23268 32508
rect 23548 32564 23604 32574
rect 23996 32564 24052 32574
rect 23548 32562 24052 32564
rect 23548 32510 23550 32562
rect 23602 32510 23998 32562
rect 24050 32510 24052 32562
rect 23548 32508 24052 32510
rect 23548 32498 23604 32508
rect 22764 32228 22820 32238
rect 22428 31164 22596 31220
rect 22652 32004 22708 32014
rect 22204 30034 22260 30044
rect 22316 30660 22372 30670
rect 22092 29934 22094 29986
rect 22146 29934 22148 29986
rect 22092 29876 22148 29934
rect 22092 29810 22148 29820
rect 21644 29586 21700 29596
rect 21756 28756 21812 28766
rect 21420 28754 21812 28756
rect 21420 28702 21422 28754
rect 21474 28702 21758 28754
rect 21810 28702 21812 28754
rect 21420 28700 21812 28702
rect 19628 28354 19684 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19516 27806 19518 27858
rect 19570 27806 19572 27858
rect 19516 27794 19572 27806
rect 21196 27860 21252 27870
rect 19404 27076 19460 27086
rect 19404 26982 19460 27020
rect 21196 27074 21252 27804
rect 21196 27022 21198 27074
rect 21250 27022 21252 27074
rect 21196 27010 21252 27022
rect 21420 26908 21476 28700
rect 21756 28690 21812 28700
rect 21868 28418 21924 28430
rect 21868 28366 21870 28418
rect 21922 28366 21924 28418
rect 21756 28084 21812 28094
rect 21868 28084 21924 28366
rect 21756 28082 21924 28084
rect 21756 28030 21758 28082
rect 21810 28030 21924 28082
rect 21756 28028 21924 28030
rect 21756 28018 21812 28028
rect 21980 27636 22036 27646
rect 21868 27580 21980 27636
rect 21868 27074 21924 27580
rect 21980 27570 22036 27580
rect 21868 27022 21870 27074
rect 21922 27022 21924 27074
rect 21868 27010 21924 27022
rect 19292 26852 19348 26862
rect 19180 26796 19292 26852
rect 18956 26786 19012 26796
rect 19068 26178 19124 26796
rect 19292 26786 19348 26796
rect 20860 26852 21476 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19964 26292 20020 26302
rect 19068 26126 19070 26178
rect 19122 26126 19124 26178
rect 19068 26114 19124 26126
rect 19292 26290 20020 26292
rect 19292 26238 19966 26290
rect 20018 26238 20020 26290
rect 19292 26236 20020 26238
rect 19292 26178 19348 26236
rect 19292 26126 19294 26178
rect 19346 26126 19348 26178
rect 18844 25666 18900 25676
rect 18788 25116 19236 25172
rect 18732 25106 18788 25116
rect 18732 24948 18788 24958
rect 18732 24854 18788 24892
rect 18844 24948 18900 24958
rect 19068 24948 19124 24958
rect 18844 24946 19068 24948
rect 18844 24894 18846 24946
rect 18898 24894 19068 24946
rect 18844 24892 19068 24894
rect 18844 24882 18900 24892
rect 19068 24882 19124 24892
rect 18620 24724 18676 24734
rect 18620 24630 18676 24668
rect 18732 23828 18788 23838
rect 18508 23772 18676 23828
rect 18396 23714 18452 23726
rect 18396 23662 18398 23714
rect 18450 23662 18452 23714
rect 18396 23604 18452 23662
rect 18620 23716 18676 23772
rect 18732 23734 18788 23772
rect 18620 23650 18676 23660
rect 18396 23548 18564 23604
rect 18396 23380 18452 23390
rect 18396 23156 18452 23324
rect 18508 23156 18564 23548
rect 18508 23100 18788 23156
rect 18396 23090 18452 23100
rect 18620 22258 18676 22270
rect 18620 22206 18622 22258
rect 18674 22206 18676 22258
rect 17724 21362 17780 21374
rect 17724 21310 17726 21362
rect 17778 21310 17780 21362
rect 17612 21252 17668 21262
rect 17276 20748 17556 20804
rect 17052 20710 17108 20748
rect 17164 20692 17220 20702
rect 17164 20690 17444 20692
rect 17164 20638 17166 20690
rect 17218 20638 17444 20690
rect 17164 20636 17444 20638
rect 17164 20626 17220 20636
rect 16716 19740 16996 19796
rect 17052 20244 17108 20254
rect 16716 19234 16772 19740
rect 16716 19182 16718 19234
rect 16770 19182 16772 19234
rect 15932 18674 16436 18676
rect 15932 18622 15934 18674
rect 15986 18622 16436 18674
rect 15932 18620 16436 18622
rect 16492 19010 16548 19022
rect 16492 18958 16494 19010
rect 16546 18958 16548 19010
rect 15932 18610 15988 18620
rect 15820 18510 15822 18562
rect 15874 18510 15876 18562
rect 15820 18498 15876 18510
rect 16268 18452 16324 18462
rect 16268 18358 16324 18396
rect 16492 18452 16548 18958
rect 16716 19012 16772 19182
rect 16828 19236 16884 19246
rect 16828 19142 16884 19180
rect 16940 19236 16996 19246
rect 17052 19236 17108 20188
rect 17388 20018 17444 20636
rect 17388 19966 17390 20018
rect 17442 19966 17444 20018
rect 17388 19954 17444 19966
rect 16940 19234 17108 19236
rect 16940 19182 16942 19234
rect 16994 19182 17108 19234
rect 16940 19180 17108 19182
rect 17164 19234 17220 19246
rect 17164 19182 17166 19234
rect 17218 19182 17220 19234
rect 16940 19170 16996 19180
rect 16716 18956 17108 19012
rect 16492 18386 16548 18396
rect 16380 18340 16436 18350
rect 16380 17892 16436 18284
rect 16828 18340 16884 18350
rect 16828 18246 16884 18284
rect 16268 17780 16324 17790
rect 16380 17780 16436 17836
rect 16268 17778 16436 17780
rect 16268 17726 16270 17778
rect 16322 17726 16436 17778
rect 16268 17724 16436 17726
rect 16604 17780 16660 17790
rect 16268 17714 16324 17724
rect 16604 17686 16660 17724
rect 17052 17778 17108 18956
rect 17052 17726 17054 17778
rect 17106 17726 17108 17778
rect 17052 17332 17108 17726
rect 17164 17780 17220 19182
rect 17164 17714 17220 17724
rect 17500 17890 17556 20748
rect 17612 20802 17668 21196
rect 17612 20750 17614 20802
rect 17666 20750 17668 20802
rect 17612 20738 17668 20750
rect 17724 20804 17780 21310
rect 17724 20738 17780 20748
rect 17724 20578 17780 20590
rect 17724 20526 17726 20578
rect 17778 20526 17780 20578
rect 17724 20468 17780 20526
rect 17836 20580 17892 20590
rect 17836 20486 17892 20524
rect 17948 20578 18004 21644
rect 18172 21644 18340 21700
rect 18396 22146 18452 22158
rect 18396 22094 18398 22146
rect 18450 22094 18452 22146
rect 18060 21028 18116 21038
rect 18060 20802 18116 20972
rect 18060 20750 18062 20802
rect 18114 20750 18116 20802
rect 18060 20738 18116 20750
rect 17948 20526 17950 20578
rect 18002 20526 18004 20578
rect 17724 20402 17780 20412
rect 17948 20468 18004 20526
rect 17948 20402 18004 20412
rect 17836 20356 17892 20366
rect 17724 20244 17780 20254
rect 17724 20150 17780 20188
rect 17836 20242 17892 20300
rect 17836 20190 17838 20242
rect 17890 20190 17892 20242
rect 17836 20178 17892 20190
rect 18060 20132 18116 20142
rect 18172 20132 18228 21644
rect 18284 21476 18340 21514
rect 18284 21410 18340 21420
rect 17948 20130 18228 20132
rect 17948 20078 18062 20130
rect 18114 20078 18228 20130
rect 17948 20076 18228 20078
rect 18284 21252 18340 21262
rect 17612 20020 17668 20030
rect 17612 20018 17892 20020
rect 17612 19966 17614 20018
rect 17666 19966 17892 20018
rect 17612 19964 17892 19966
rect 17612 19954 17668 19964
rect 17836 19908 17892 19964
rect 17724 19236 17780 19246
rect 17724 19142 17780 19180
rect 17724 19012 17780 19022
rect 17836 19012 17892 19852
rect 17780 18956 17892 19012
rect 17724 18674 17780 18956
rect 17724 18622 17726 18674
rect 17778 18622 17780 18674
rect 17724 18610 17780 18622
rect 17836 18452 17892 18462
rect 17836 18358 17892 18396
rect 17500 17838 17502 17890
rect 17554 17838 17556 17890
rect 17500 17444 17556 17838
rect 17948 17780 18004 20076
rect 18060 20066 18116 20076
rect 18284 18900 18340 21196
rect 18396 20916 18452 22094
rect 18396 20850 18452 20860
rect 18508 21588 18564 21598
rect 18396 20468 18452 20478
rect 18396 20132 18452 20412
rect 18508 20244 18564 21532
rect 18620 21140 18676 22206
rect 18732 22146 18788 23100
rect 18732 22094 18734 22146
rect 18786 22094 18788 22146
rect 18732 22036 18788 22094
rect 18956 22148 19012 22158
rect 18956 22054 19012 22092
rect 18732 21970 18788 21980
rect 18620 21074 18676 21084
rect 19068 21028 19124 21038
rect 18732 21026 19124 21028
rect 18732 20974 19070 21026
rect 19122 20974 19124 21026
rect 18732 20972 19124 20974
rect 18620 20914 18676 20926
rect 18620 20862 18622 20914
rect 18674 20862 18676 20914
rect 18620 20804 18676 20862
rect 18620 20738 18676 20748
rect 18620 20580 18676 20590
rect 18732 20580 18788 20972
rect 19068 20962 19124 20972
rect 18844 20692 18900 20702
rect 18844 20598 18900 20636
rect 18620 20578 18788 20580
rect 18620 20526 18622 20578
rect 18674 20526 18788 20578
rect 18620 20524 18788 20526
rect 18620 20514 18676 20524
rect 18620 20244 18676 20254
rect 18508 20242 18676 20244
rect 18508 20190 18622 20242
rect 18674 20190 18676 20242
rect 18508 20188 18676 20190
rect 18620 20178 18676 20188
rect 18396 20076 18564 20132
rect 18060 18844 18340 18900
rect 18060 18674 18116 18844
rect 18060 18622 18062 18674
rect 18114 18622 18116 18674
rect 18060 18340 18116 18622
rect 18508 18676 18564 20076
rect 18732 20020 18788 20524
rect 18732 19954 18788 19964
rect 19180 19906 19236 25116
rect 19292 25060 19348 26126
rect 19964 26180 20020 26236
rect 19964 26114 20020 26124
rect 20860 26292 20916 26852
rect 22316 26740 22372 30604
rect 22316 26674 22372 26684
rect 22428 26516 22484 31164
rect 22540 30884 22596 30894
rect 22652 30884 22708 31948
rect 22764 31554 22820 32172
rect 23436 31780 23492 31790
rect 23436 31686 23492 31724
rect 23212 31668 23268 31678
rect 23212 31574 23268 31612
rect 22764 31502 22766 31554
rect 22818 31502 22820 31554
rect 22764 31490 22820 31502
rect 23324 31556 23380 31566
rect 23772 31556 23828 32508
rect 23996 32498 24052 32508
rect 24220 32562 24276 32574
rect 24220 32510 24222 32562
rect 24274 32510 24276 32562
rect 24108 32228 24164 32238
rect 24220 32228 24276 32510
rect 24164 32172 24276 32228
rect 24668 32564 24724 32574
rect 24780 32564 24836 33070
rect 24668 32562 24836 32564
rect 24668 32510 24670 32562
rect 24722 32510 24836 32562
rect 24668 32508 24836 32510
rect 24108 32162 24164 32172
rect 24220 31892 24276 31902
rect 23884 31890 24276 31892
rect 23884 31838 24222 31890
rect 24274 31838 24276 31890
rect 23884 31836 24276 31838
rect 23884 31778 23940 31836
rect 24220 31826 24276 31836
rect 24668 31892 24724 32508
rect 24668 31826 24724 31836
rect 23884 31726 23886 31778
rect 23938 31726 23940 31778
rect 23884 31714 23940 31726
rect 24444 31780 24500 31790
rect 24444 31686 24500 31724
rect 24108 31666 24164 31678
rect 24108 31614 24110 31666
rect 24162 31614 24164 31666
rect 24108 31556 24164 31614
rect 23772 31500 24164 31556
rect 23324 31462 23380 31500
rect 22876 30994 22932 31006
rect 22876 30942 22878 30994
rect 22930 30942 22932 30994
rect 22876 30884 22932 30942
rect 22540 30882 22932 30884
rect 22540 30830 22542 30882
rect 22594 30830 22932 30882
rect 22540 30828 22932 30830
rect 22540 30818 22596 30828
rect 22764 30212 22820 30222
rect 22876 30212 22932 30828
rect 23324 30882 23380 30894
rect 23324 30830 23326 30882
rect 23378 30830 23380 30882
rect 23324 30660 23380 30830
rect 23324 30594 23380 30604
rect 23324 30212 23380 30222
rect 25564 30212 25620 35868
rect 25676 35922 25732 37212
rect 25676 35870 25678 35922
rect 25730 35870 25732 35922
rect 25676 35858 25732 35870
rect 25788 35588 25844 37324
rect 25900 37268 25956 37278
rect 25900 36932 25956 37212
rect 25900 36866 25956 36876
rect 26572 37266 26628 37278
rect 26572 37214 26574 37266
rect 26626 37214 26628 37266
rect 26236 36820 26292 36830
rect 25788 35522 25844 35532
rect 26124 36372 26180 36382
rect 26124 35138 26180 36316
rect 26236 35922 26292 36764
rect 26572 36596 26628 37214
rect 26572 36530 26628 36540
rect 26236 35870 26238 35922
rect 26290 35870 26292 35922
rect 26236 35858 26292 35870
rect 26572 36258 26628 36270
rect 26572 36206 26574 36258
rect 26626 36206 26628 36258
rect 26572 35922 26628 36206
rect 26572 35870 26574 35922
rect 26626 35870 26628 35922
rect 26572 35858 26628 35870
rect 26684 35700 26740 35710
rect 26684 35606 26740 35644
rect 26908 35476 26964 38556
rect 27020 38546 27076 38556
rect 27132 36036 27188 38780
rect 27244 38050 27300 38062
rect 27244 37998 27246 38050
rect 27298 37998 27300 38050
rect 27244 37044 27300 37998
rect 27580 37492 27636 41200
rect 28476 38610 28532 38622
rect 28476 38558 28478 38610
rect 28530 38558 28532 38610
rect 28476 38050 28532 38558
rect 28812 38612 28868 38622
rect 28812 38162 28868 38556
rect 28924 38276 28980 41200
rect 31612 38668 31668 41200
rect 32284 39508 32340 41200
rect 32284 39452 32788 39508
rect 31612 38612 31892 38668
rect 28924 38210 28980 38220
rect 30380 38276 30436 38286
rect 28812 38110 28814 38162
rect 28866 38110 28868 38162
rect 28812 38098 28868 38110
rect 30380 38162 30436 38220
rect 30380 38110 30382 38162
rect 30434 38110 30436 38162
rect 30380 38098 30436 38110
rect 28476 37998 28478 38050
rect 28530 37998 28532 38050
rect 28476 37986 28532 37998
rect 27804 37828 27860 37838
rect 29708 37828 29764 37838
rect 29932 37828 29988 37838
rect 27804 37734 27860 37772
rect 29484 37826 29764 37828
rect 29484 37774 29710 37826
rect 29762 37774 29764 37826
rect 29484 37772 29764 37774
rect 27580 37426 27636 37436
rect 28924 37490 28980 37502
rect 28924 37438 28926 37490
rect 28978 37438 28980 37490
rect 28700 37380 28756 37390
rect 27916 37268 27972 37278
rect 27244 36706 27300 36988
rect 27244 36654 27246 36706
rect 27298 36654 27300 36706
rect 27244 36642 27300 36654
rect 27804 37212 27916 37268
rect 27580 36596 27636 36606
rect 27580 36502 27636 36540
rect 27468 36372 27524 36382
rect 27692 36372 27748 36382
rect 27468 36370 27636 36372
rect 27468 36318 27470 36370
rect 27522 36318 27636 36370
rect 27468 36316 27636 36318
rect 27468 36306 27524 36316
rect 27132 35980 27412 36036
rect 27356 35924 27412 35980
rect 27132 35812 27188 35822
rect 26124 35086 26126 35138
rect 26178 35086 26180 35138
rect 25676 34916 25732 34926
rect 25676 34822 25732 34860
rect 26124 34690 26180 35086
rect 26684 35420 26964 35476
rect 27020 35810 27188 35812
rect 27020 35758 27134 35810
rect 27186 35758 27188 35810
rect 27020 35756 27188 35758
rect 26572 34804 26628 34814
rect 26572 34710 26628 34748
rect 26124 34638 26126 34690
rect 26178 34638 26180 34690
rect 26124 34580 26180 34638
rect 26124 34524 26404 34580
rect 25676 34244 25732 34254
rect 25676 34150 25732 34188
rect 26236 34132 26292 34142
rect 26236 34038 26292 34076
rect 26124 34020 26180 34030
rect 26124 33926 26180 33964
rect 26124 33572 26180 33582
rect 26124 33458 26180 33516
rect 26124 33406 26126 33458
rect 26178 33406 26180 33458
rect 26124 33394 26180 33406
rect 26236 33124 26292 33134
rect 26236 33030 26292 33068
rect 26348 32452 26404 34524
rect 26460 34020 26516 34030
rect 26460 33684 26516 33964
rect 26460 33618 26516 33628
rect 26236 32396 26404 32452
rect 25676 31780 25732 31790
rect 25676 31686 25732 31724
rect 26012 31668 26068 31678
rect 26012 31574 26068 31612
rect 22764 30210 23380 30212
rect 22764 30158 22766 30210
rect 22818 30158 23326 30210
rect 23378 30158 23380 30210
rect 22764 30156 23380 30158
rect 22764 30146 22820 30156
rect 22540 29652 22596 29662
rect 22540 28082 22596 29596
rect 22540 28030 22542 28082
rect 22594 28030 22596 28082
rect 22540 28018 22596 28030
rect 22652 28644 22708 28654
rect 22988 28644 23044 28654
rect 22652 28642 23044 28644
rect 22652 28590 22654 28642
rect 22706 28590 22990 28642
rect 23042 28590 23044 28642
rect 22652 28588 23044 28590
rect 22652 27860 22708 28588
rect 22988 28578 23044 28588
rect 22764 28084 22820 28094
rect 22764 28082 23156 28084
rect 22764 28030 22766 28082
rect 22818 28030 23156 28082
rect 22764 28028 23156 28030
rect 22764 28018 22820 28028
rect 22652 27794 22708 27804
rect 22988 27858 23044 27870
rect 22988 27806 22990 27858
rect 23042 27806 23044 27858
rect 22876 27746 22932 27758
rect 22876 27694 22878 27746
rect 22930 27694 22932 27746
rect 22876 27636 22932 27694
rect 22876 27570 22932 27580
rect 22988 27748 23044 27806
rect 22988 26908 23044 27692
rect 19404 26068 19460 26078
rect 19404 26066 19572 26068
rect 19404 26014 19406 26066
rect 19458 26014 19572 26066
rect 19404 26012 19572 26014
rect 19404 26002 19460 26012
rect 19516 25394 19572 26012
rect 19516 25342 19518 25394
rect 19570 25342 19572 25394
rect 19516 25330 19572 25342
rect 19628 25732 19684 25742
rect 19292 24994 19348 25004
rect 19516 24948 19572 24958
rect 19404 24834 19460 24846
rect 19404 24782 19406 24834
rect 19458 24782 19460 24834
rect 19292 24724 19348 24734
rect 19404 24724 19460 24782
rect 19292 24722 19460 24724
rect 19292 24670 19294 24722
rect 19346 24670 19460 24722
rect 19292 24668 19460 24670
rect 19292 24658 19348 24668
rect 19404 24052 19460 24062
rect 19516 24052 19572 24892
rect 19628 24946 19684 25676
rect 20300 25732 20356 25742
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20300 24948 20356 25676
rect 20636 25396 20692 25406
rect 20636 25284 20692 25340
rect 19628 24894 19630 24946
rect 19682 24894 19684 24946
rect 19628 24882 19684 24894
rect 20076 24946 20356 24948
rect 20076 24894 20302 24946
rect 20354 24894 20356 24946
rect 20076 24892 20356 24894
rect 19740 24836 19796 24846
rect 19740 24612 19796 24780
rect 19740 24546 19796 24556
rect 19292 24050 19572 24052
rect 19292 23998 19406 24050
rect 19458 23998 19572 24050
rect 19292 23996 19572 23998
rect 19292 23380 19348 23996
rect 19404 23986 19460 23996
rect 20076 23938 20132 24892
rect 20300 24882 20356 24892
rect 20412 25282 20692 25284
rect 20412 25230 20638 25282
rect 20690 25230 20692 25282
rect 20412 25228 20692 25230
rect 20076 23886 20078 23938
rect 20130 23886 20132 23938
rect 20076 23874 20132 23886
rect 20188 24722 20244 24734
rect 20188 24670 20190 24722
rect 20242 24670 20244 24722
rect 20188 24052 20244 24670
rect 20300 24612 20356 24622
rect 20412 24612 20468 25228
rect 20636 25218 20692 25228
rect 20860 25060 20916 26236
rect 21868 26460 22484 26516
rect 22652 26852 23044 26908
rect 21532 26178 21588 26190
rect 21532 26126 21534 26178
rect 21586 26126 21588 26178
rect 21532 25730 21588 26126
rect 21532 25678 21534 25730
rect 21586 25678 21588 25730
rect 21532 25666 21588 25678
rect 20636 25004 20916 25060
rect 21420 25394 21476 25406
rect 21420 25342 21422 25394
rect 21474 25342 21476 25394
rect 20524 24836 20580 24846
rect 20524 24742 20580 24780
rect 20636 24612 20692 25004
rect 21196 24948 21252 24958
rect 21420 24948 21476 25342
rect 20860 24946 21476 24948
rect 20860 24894 21198 24946
rect 21250 24894 21476 24946
rect 20860 24892 21476 24894
rect 21532 25282 21588 25294
rect 21532 25230 21534 25282
rect 21586 25230 21588 25282
rect 20356 24556 20468 24612
rect 20524 24556 20692 24612
rect 20748 24722 20804 24734
rect 20748 24670 20750 24722
rect 20802 24670 20804 24722
rect 20300 24546 20356 24556
rect 20300 24052 20356 24062
rect 20188 24050 20356 24052
rect 20188 23998 20302 24050
rect 20354 23998 20356 24050
rect 20188 23996 20356 23998
rect 19516 23828 19572 23838
rect 19292 23314 19348 23324
rect 19404 23716 19460 23726
rect 19292 23044 19348 23054
rect 19292 22950 19348 22988
rect 19292 22146 19348 22158
rect 19292 22094 19294 22146
rect 19346 22094 19348 22146
rect 19292 22036 19348 22094
rect 19292 21970 19348 21980
rect 19292 21812 19348 21822
rect 19292 20914 19348 21756
rect 19292 20862 19294 20914
rect 19346 20862 19348 20914
rect 19292 20850 19348 20862
rect 19180 19854 19182 19906
rect 19234 19854 19236 19906
rect 19180 19842 19236 19854
rect 18732 18676 18788 18686
rect 18508 18674 18788 18676
rect 18508 18622 18734 18674
rect 18786 18622 18788 18674
rect 18508 18620 18788 18622
rect 18732 18610 18788 18620
rect 19180 18564 19236 18574
rect 18060 18274 18116 18284
rect 18172 18450 18228 18462
rect 18172 18398 18174 18450
rect 18226 18398 18228 18450
rect 18172 17890 18228 18398
rect 19180 18450 19236 18508
rect 19180 18398 19182 18450
rect 19234 18398 19236 18450
rect 19180 18386 19236 18398
rect 19404 18228 19460 23660
rect 19516 19124 19572 23772
rect 19836 23548 20100 23558
rect 19628 23492 19684 23502
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 23378 19684 23436
rect 19628 23326 19630 23378
rect 19682 23326 19684 23378
rect 19628 23268 19684 23326
rect 19628 23202 19684 23212
rect 19964 23380 20020 23390
rect 19964 23044 20020 23324
rect 20076 23380 20132 23390
rect 20188 23380 20244 23996
rect 20300 23986 20356 23996
rect 20076 23378 20244 23380
rect 20076 23326 20078 23378
rect 20130 23326 20244 23378
rect 20076 23324 20244 23326
rect 20076 23314 20132 23324
rect 20412 23268 20468 23278
rect 20412 23156 20468 23212
rect 19740 22148 19796 22158
rect 19628 22146 19796 22148
rect 19628 22094 19742 22146
rect 19794 22094 19796 22146
rect 19628 22092 19796 22094
rect 19628 21026 19684 22092
rect 19740 22082 19796 22092
rect 19964 22148 20020 22988
rect 19964 22082 20020 22092
rect 20188 23154 20468 23156
rect 20188 23102 20414 23154
rect 20466 23102 20468 23154
rect 20188 23100 20468 23102
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19628 20974 19630 21026
rect 19682 20974 19684 21026
rect 19628 20962 19684 20974
rect 19852 21252 19908 21262
rect 19852 20692 19908 21196
rect 20188 21140 20244 23100
rect 20412 23090 20468 23100
rect 20524 22932 20580 24556
rect 20636 23940 20692 23950
rect 20636 23548 20692 23884
rect 20748 23828 20804 24670
rect 20748 23734 20804 23772
rect 20636 23492 20804 23548
rect 20748 23380 20804 23492
rect 20748 23314 20804 23324
rect 20636 23156 20692 23166
rect 20860 23156 20916 24892
rect 21196 24882 21252 24892
rect 21532 24836 21588 25230
rect 21868 24948 21924 26460
rect 22540 26404 22596 26414
rect 22428 26348 22540 26404
rect 21980 26290 22036 26302
rect 21980 26238 21982 26290
rect 22034 26238 22036 26290
rect 21980 25172 22036 26238
rect 22428 26290 22484 26348
rect 22540 26338 22596 26348
rect 22428 26238 22430 26290
rect 22482 26238 22484 26290
rect 22428 26226 22484 26238
rect 22428 25508 22484 25518
rect 21980 25106 22036 25116
rect 22092 25506 22484 25508
rect 22092 25454 22430 25506
rect 22482 25454 22484 25506
rect 22092 25452 22484 25454
rect 21868 24892 22036 24948
rect 21532 24770 21588 24780
rect 21084 24724 21140 24734
rect 20972 24722 21140 24724
rect 20972 24670 21086 24722
rect 21138 24670 21140 24722
rect 20972 24668 21140 24670
rect 20972 23940 21028 24668
rect 21084 24658 21140 24668
rect 21308 24724 21364 24734
rect 21644 24724 21700 24734
rect 21308 24722 21476 24724
rect 21308 24670 21310 24722
rect 21362 24670 21476 24722
rect 21308 24668 21476 24670
rect 21308 24658 21364 24668
rect 21420 23940 21476 24668
rect 21700 24668 21812 24724
rect 21644 24658 21700 24668
rect 21756 24050 21812 24668
rect 21756 23998 21758 24050
rect 21810 23998 21812 24050
rect 21756 23986 21812 23998
rect 21644 23940 21700 23950
rect 21420 23884 21644 23940
rect 20972 23874 21028 23884
rect 21308 23826 21364 23838
rect 21308 23774 21310 23826
rect 21362 23774 21364 23826
rect 21308 23604 21364 23774
rect 21532 23716 21588 23726
rect 20972 23548 21364 23604
rect 21420 23714 21588 23716
rect 21420 23662 21534 23714
rect 21586 23662 21588 23714
rect 21420 23660 21588 23662
rect 20972 23378 21028 23548
rect 21420 23492 21476 23660
rect 21532 23650 21588 23660
rect 21644 23492 21700 23884
rect 21196 23436 21476 23492
rect 21532 23436 21700 23492
rect 21756 23714 21812 23726
rect 21756 23662 21758 23714
rect 21810 23662 21812 23714
rect 20972 23326 20974 23378
rect 21026 23326 21028 23378
rect 20972 23314 21028 23326
rect 21084 23380 21140 23390
rect 20636 23154 20916 23156
rect 20636 23102 20638 23154
rect 20690 23102 20916 23154
rect 20636 23100 20916 23102
rect 20972 23156 21028 23166
rect 20636 23090 20692 23100
rect 20412 22876 20580 22932
rect 20300 22146 20356 22158
rect 20300 22094 20302 22146
rect 20354 22094 20356 22146
rect 20300 22036 20356 22094
rect 20300 21970 20356 21980
rect 20412 21364 20468 22876
rect 20972 22372 21028 23100
rect 21084 23044 21140 23324
rect 21196 23378 21252 23436
rect 21196 23326 21198 23378
rect 21250 23326 21252 23378
rect 21196 23314 21252 23326
rect 21196 23044 21252 23054
rect 21084 22988 21196 23044
rect 21196 22978 21252 22988
rect 21532 22820 21588 23436
rect 21756 23268 21812 23662
rect 21868 23714 21924 23726
rect 21868 23662 21870 23714
rect 21922 23662 21924 23714
rect 21868 23380 21924 23662
rect 21980 23492 22036 24892
rect 22092 24724 22148 25452
rect 22428 25442 22484 25452
rect 22540 25284 22596 25294
rect 22428 25172 22484 25182
rect 22092 24630 22148 24668
rect 22316 25116 22428 25172
rect 22204 24610 22260 24622
rect 22204 24558 22206 24610
rect 22258 24558 22260 24610
rect 21980 23426 22036 23436
rect 22092 23828 22148 23838
rect 21868 23314 21924 23324
rect 21644 23212 21812 23268
rect 21644 23156 21700 23212
rect 22092 23210 22148 23772
rect 22092 23158 22094 23210
rect 22146 23158 22148 23210
rect 22092 23146 22148 23158
rect 21644 23090 21700 23100
rect 21868 23044 21924 23054
rect 21868 22950 21924 22988
rect 21644 22930 21700 22942
rect 21644 22878 21646 22930
rect 21698 22878 21700 22930
rect 21644 22820 21700 22878
rect 20636 22316 21028 22372
rect 21420 22764 21700 22820
rect 21756 22820 21812 22830
rect 19852 20598 19908 20636
rect 20076 21084 20244 21140
rect 20300 21308 20468 21364
rect 20524 22148 20580 22158
rect 20076 20580 20132 21084
rect 20188 20916 20244 20926
rect 20188 20822 20244 20860
rect 20076 20524 20244 20580
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19516 19058 19572 19068
rect 19852 20018 19908 20030
rect 19852 19966 19854 20018
rect 19906 19966 19908 20018
rect 19852 19012 19908 19966
rect 19628 18956 19908 19012
rect 19628 18452 19684 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19740 18452 19796 18462
rect 19628 18450 19796 18452
rect 19628 18398 19742 18450
rect 19794 18398 19796 18450
rect 19628 18396 19796 18398
rect 19404 18162 19460 18172
rect 18172 17838 18174 17890
rect 18226 17838 18228 17890
rect 18060 17780 18116 17790
rect 17948 17778 18116 17780
rect 17948 17726 18062 17778
rect 18114 17726 18116 17778
rect 17948 17724 18116 17726
rect 18060 17714 18116 17724
rect 18172 17668 18228 17838
rect 18956 18116 19012 18126
rect 18396 17780 18452 17790
rect 18396 17686 18452 17724
rect 18956 17778 19012 18060
rect 19740 17892 19796 18396
rect 20188 18340 20244 20524
rect 20300 19348 20356 21308
rect 20524 20916 20580 22092
rect 20636 21026 20692 22316
rect 20748 22148 20804 22158
rect 20748 22054 20804 22092
rect 21420 21812 21476 22764
rect 21644 22484 21700 22494
rect 21756 22484 21812 22764
rect 21644 22482 21812 22484
rect 21644 22430 21646 22482
rect 21698 22430 21812 22482
rect 21644 22428 21812 22430
rect 21868 22596 21924 22606
rect 21644 22418 21700 22428
rect 21756 22260 21812 22270
rect 21868 22260 21924 22540
rect 22204 22596 22260 24558
rect 22316 23156 22372 25116
rect 22428 25106 22484 25116
rect 22428 23940 22484 23950
rect 22428 23846 22484 23884
rect 22428 23156 22484 23166
rect 22316 23154 22484 23156
rect 22316 23102 22430 23154
rect 22482 23102 22484 23154
rect 22316 23100 22484 23102
rect 22428 23090 22484 23100
rect 22204 22482 22260 22540
rect 22204 22430 22206 22482
rect 22258 22430 22260 22482
rect 22204 22418 22260 22430
rect 21756 22258 21924 22260
rect 21756 22206 21758 22258
rect 21810 22206 21924 22258
rect 21756 22204 21924 22206
rect 22428 22258 22484 22270
rect 22428 22206 22430 22258
rect 22482 22206 22484 22258
rect 21756 22194 21812 22204
rect 21420 21746 21476 21756
rect 21532 22146 21588 22158
rect 21532 22094 21534 22146
rect 21586 22094 21588 22146
rect 21532 22036 21588 22094
rect 20636 20974 20638 21026
rect 20690 20974 20692 21026
rect 20636 20962 20692 20974
rect 20748 21700 20804 21710
rect 20524 20692 20580 20860
rect 20748 20802 20804 21644
rect 20748 20750 20750 20802
rect 20802 20750 20804 20802
rect 20748 20738 20804 20750
rect 20636 20692 20692 20702
rect 20524 20690 20692 20692
rect 20524 20638 20638 20690
rect 20690 20638 20692 20690
rect 20524 20636 20692 20638
rect 20636 20626 20692 20636
rect 20860 20692 20916 20702
rect 20524 20018 20580 20030
rect 20524 19966 20526 20018
rect 20578 19966 20580 20018
rect 20412 19348 20468 19358
rect 20300 19292 20412 19348
rect 20412 19282 20468 19292
rect 20300 19012 20356 19022
rect 20300 18918 20356 18956
rect 19740 17826 19796 17836
rect 19852 18284 20244 18340
rect 20412 18338 20468 18350
rect 20412 18286 20414 18338
rect 20466 18286 20468 18338
rect 18956 17726 18958 17778
rect 19010 17726 19012 17778
rect 18956 17714 19012 17726
rect 19292 17780 19348 17790
rect 18172 17602 18228 17612
rect 17052 17266 17108 17276
rect 17388 17442 17556 17444
rect 17388 17390 17502 17442
rect 17554 17390 17556 17442
rect 17388 17388 17556 17390
rect 15484 17054 15486 17106
rect 15538 17054 15540 17106
rect 15484 17042 15540 17054
rect 14812 16996 14868 17006
rect 14812 16902 14868 16940
rect 17388 16996 17444 17388
rect 17500 17378 17556 17388
rect 19292 17106 19348 17724
rect 19852 17780 19908 18284
rect 20412 18228 20468 18286
rect 20412 18162 20468 18172
rect 19852 17666 19908 17724
rect 19964 18116 20020 18126
rect 19964 17778 20020 18060
rect 20412 17892 20468 17902
rect 20412 17798 20468 17836
rect 19964 17726 19966 17778
rect 20018 17726 20020 17778
rect 19964 17714 20020 17726
rect 19852 17614 19854 17666
rect 19906 17614 19908 17666
rect 19852 17602 19908 17614
rect 20300 17668 20356 17678
rect 20300 17666 20468 17668
rect 20300 17614 20302 17666
rect 20354 17614 20468 17666
rect 20300 17612 20468 17614
rect 20300 17602 20356 17612
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19292 17054 19294 17106
rect 19346 17054 19348 17106
rect 19292 17042 19348 17054
rect 17388 16930 17444 16940
rect 17500 16994 17556 17006
rect 17500 16942 17502 16994
rect 17554 16942 17556 16994
rect 15260 16882 15316 16894
rect 15260 16830 15262 16882
rect 15314 16830 15316 16882
rect 15260 16772 15316 16830
rect 15932 16884 15988 16894
rect 15932 16790 15988 16828
rect 17276 16884 17332 16894
rect 17276 16790 17332 16828
rect 15260 16706 15316 16716
rect 15372 16770 15428 16782
rect 15372 16718 15374 16770
rect 15426 16718 15428 16770
rect 15372 16436 15428 16718
rect 14252 16210 14756 16212
rect 14252 16158 14254 16210
rect 14306 16158 14756 16210
rect 14252 16156 14756 16158
rect 11116 15262 11118 15314
rect 11170 15262 11172 15314
rect 11116 15250 11172 15262
rect 14140 14644 14196 14654
rect 14252 14644 14308 16156
rect 14700 16098 14756 16156
rect 14700 16046 14702 16098
rect 14754 16046 14756 16098
rect 14700 16034 14756 16046
rect 15148 16380 15428 16436
rect 15596 16772 15652 16782
rect 15148 16098 15204 16380
rect 15148 16046 15150 16098
rect 15202 16046 15204 16098
rect 15148 16034 15204 16046
rect 14364 15540 14420 15550
rect 14364 15446 14420 15484
rect 15596 15538 15652 16716
rect 16268 16772 16324 16782
rect 16268 16678 16324 16716
rect 16828 16772 16884 16782
rect 16828 16678 16884 16716
rect 15596 15486 15598 15538
rect 15650 15486 15652 15538
rect 15596 15474 15652 15486
rect 15820 16548 15876 16558
rect 15820 15538 15876 16492
rect 17500 16324 17556 16942
rect 18396 16994 18452 17006
rect 18396 16942 18398 16994
rect 18450 16942 18452 16994
rect 17500 16258 17556 16268
rect 17612 16882 17668 16894
rect 17612 16830 17614 16882
rect 17666 16830 17668 16882
rect 17612 16772 17668 16830
rect 17388 15876 17444 15886
rect 15820 15486 15822 15538
rect 15874 15486 15876 15538
rect 15820 15474 15876 15486
rect 16828 15874 17444 15876
rect 16828 15822 17390 15874
rect 17442 15822 17444 15874
rect 16828 15820 17444 15822
rect 16828 15538 16884 15820
rect 17388 15810 17444 15820
rect 16828 15486 16830 15538
rect 16882 15486 16884 15538
rect 16828 15474 16884 15486
rect 17500 15540 17556 15550
rect 17500 15446 17556 15484
rect 14476 15428 14532 15438
rect 14476 15148 14532 15372
rect 17612 15426 17668 16716
rect 18284 16882 18340 16894
rect 18284 16830 18286 16882
rect 18338 16830 18340 16882
rect 18172 16324 18228 16334
rect 18172 16230 18228 16268
rect 18284 16100 18340 16830
rect 18396 16772 18452 16942
rect 19964 16884 20020 16894
rect 18452 16716 18564 16772
rect 18396 16706 18452 16716
rect 18396 16100 18452 16110
rect 18284 16044 18396 16100
rect 17612 15374 17614 15426
rect 17666 15374 17668 15426
rect 16268 15316 16324 15326
rect 15372 15204 15428 15242
rect 16268 15222 16324 15260
rect 17276 15316 17332 15326
rect 15708 15202 15764 15214
rect 15708 15150 15710 15202
rect 15762 15150 15764 15202
rect 15708 15148 15764 15150
rect 14476 15092 14756 15148
rect 15372 15138 15428 15148
rect 14140 14642 14308 14644
rect 14140 14590 14142 14642
rect 14194 14590 14308 14642
rect 14140 14588 14308 14590
rect 14140 14578 14196 14588
rect 10668 14466 10724 14476
rect 13692 14532 13748 14542
rect 9660 13634 10052 13636
rect 9660 13582 9662 13634
rect 9714 13582 10052 13634
rect 9660 13580 10052 13582
rect 9660 13570 9716 13580
rect 7308 13094 7364 13132
rect 7420 13186 8148 13188
rect 7420 13134 7534 13186
rect 7586 13134 8148 13186
rect 7420 13132 8148 13134
rect 6524 13022 6526 13074
rect 6578 13022 6580 13074
rect 6524 13010 6580 13022
rect 2268 12870 2324 12908
rect 4844 12964 4900 12974
rect 6076 12964 6132 12974
rect 4844 12404 4900 12908
rect 5964 12962 6132 12964
rect 5964 12910 6078 12962
rect 6130 12910 6132 12962
rect 5964 12908 6132 12910
rect 4844 12402 5236 12404
rect 4844 12350 4846 12402
rect 4898 12350 5236 12402
rect 4844 12348 5236 12350
rect 4844 12338 4900 12348
rect 5180 12178 5236 12348
rect 5180 12126 5182 12178
rect 5234 12126 5236 12178
rect 5180 12114 5236 12126
rect 5964 12066 6020 12908
rect 6076 12898 6132 12908
rect 7420 12628 7476 13132
rect 7532 13122 7588 13132
rect 7980 12964 8036 12974
rect 7980 12870 8036 12908
rect 7644 12852 7700 12862
rect 7644 12758 7700 12796
rect 5964 12014 5966 12066
rect 6018 12014 6020 12066
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 5964 11620 6020 12014
rect 6972 12572 7476 12628
rect 5964 11554 6020 11564
rect 6860 11620 6916 11630
rect 6860 11526 6916 11564
rect 6972 11506 7028 12572
rect 8092 12066 8148 13132
rect 8540 12964 8596 12974
rect 8540 12292 8596 12908
rect 8764 12852 8820 12862
rect 8764 12758 8820 12796
rect 8540 12198 8596 12236
rect 9996 12292 10052 13580
rect 13692 13858 13748 14476
rect 14252 14532 14308 14588
rect 14700 14642 14756 15092
rect 14700 14590 14702 14642
rect 14754 14590 14756 14642
rect 14700 14578 14756 14590
rect 15484 15092 15764 15148
rect 16716 15204 16772 15242
rect 17276 15222 17332 15260
rect 16716 15138 16772 15148
rect 17612 15148 17668 15374
rect 18396 15540 18452 16044
rect 18060 15204 18116 15242
rect 17612 15092 17892 15148
rect 18060 15138 18116 15148
rect 18396 15148 18452 15484
rect 18508 15426 18564 16716
rect 18732 16770 18788 16782
rect 18732 16718 18734 16770
rect 18786 16718 18788 16770
rect 18732 16436 18788 16718
rect 19628 16772 19684 16782
rect 19852 16772 19908 16782
rect 19684 16770 19908 16772
rect 19684 16718 19854 16770
rect 19906 16718 19908 16770
rect 19684 16716 19908 16718
rect 18732 16370 18788 16380
rect 19516 16436 19572 16446
rect 18508 15374 18510 15426
rect 18562 15374 18564 15426
rect 18508 15362 18564 15374
rect 18620 16324 18676 16334
rect 18620 15316 18676 16268
rect 19404 16212 19460 16222
rect 19292 16100 19348 16110
rect 19292 16006 19348 16044
rect 19180 15428 19236 15438
rect 18732 15316 18788 15326
rect 18620 15314 18788 15316
rect 18620 15262 18734 15314
rect 18786 15262 18788 15314
rect 18620 15260 18788 15262
rect 18732 15204 18788 15260
rect 14252 14466 14308 14476
rect 14924 14532 14980 14542
rect 13692 13806 13694 13858
rect 13746 13806 13748 13858
rect 10892 13076 10948 13086
rect 10892 12982 10948 13020
rect 12012 13076 12068 13086
rect 12012 12982 12068 13020
rect 12460 13076 12516 13086
rect 12908 13076 12964 13086
rect 13692 13076 13748 13806
rect 12460 13074 13748 13076
rect 12460 13022 12462 13074
rect 12514 13022 12910 13074
rect 12962 13022 13694 13074
rect 13746 13022 13748 13074
rect 12460 13020 13748 13022
rect 12460 13010 12516 13020
rect 12908 13010 12964 13020
rect 8092 12014 8094 12066
rect 8146 12014 8148 12066
rect 8092 12002 8148 12014
rect 6972 11454 6974 11506
rect 7026 11454 7028 11506
rect 6972 11442 7028 11454
rect 9436 11394 9492 11406
rect 9996 11396 10052 12236
rect 11228 12850 11284 12862
rect 11228 12798 11230 12850
rect 11282 12798 11284 12850
rect 11228 12740 11284 12798
rect 10668 12068 10724 12078
rect 10668 12066 10836 12068
rect 10668 12014 10670 12066
rect 10722 12014 10836 12066
rect 10668 12012 10836 12014
rect 10668 12002 10724 12012
rect 9436 11342 9438 11394
rect 9490 11342 9492 11394
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 9436 10052 9492 11342
rect 9772 11394 10052 11396
rect 9772 11342 9998 11394
rect 10050 11342 10052 11394
rect 9772 11340 10052 11342
rect 9660 11172 9716 11182
rect 9660 11078 9716 11116
rect 9660 10612 9716 10622
rect 9772 10612 9828 11340
rect 9996 11330 10052 11340
rect 10780 11284 10836 12012
rect 10780 11190 10836 11228
rect 10332 11172 10388 11182
rect 10332 10722 10388 11116
rect 10332 10670 10334 10722
rect 10386 10670 10388 10722
rect 10332 10658 10388 10670
rect 9660 10610 9828 10612
rect 9660 10558 9662 10610
rect 9714 10558 9828 10610
rect 9660 10556 9828 10558
rect 9660 10546 9716 10556
rect 9436 9986 9492 9996
rect 10780 10052 10836 10062
rect 10780 9958 10836 9996
rect 11116 10052 11172 10062
rect 11228 10052 11284 12684
rect 11340 12738 11396 12750
rect 11340 12686 11342 12738
rect 11394 12686 11396 12738
rect 11340 11956 11396 12686
rect 11340 11890 11396 11900
rect 11452 12738 11508 12750
rect 11452 12686 11454 12738
rect 11506 12686 11508 12738
rect 11116 10050 11284 10052
rect 11116 9998 11118 10050
rect 11170 9998 11284 10050
rect 11116 9996 11284 9998
rect 11452 10500 11508 12686
rect 11900 12740 11956 12750
rect 11900 12646 11956 12684
rect 13468 12180 13524 13020
rect 13692 13010 13748 13020
rect 14700 13076 14756 13086
rect 14364 12850 14420 12862
rect 14364 12798 14366 12850
rect 14418 12798 14420 12850
rect 13916 12180 13972 12190
rect 13468 12178 13972 12180
rect 13468 12126 13470 12178
rect 13522 12126 13918 12178
rect 13970 12126 13972 12178
rect 13468 12124 13972 12126
rect 13468 12114 13524 12124
rect 12796 12066 12852 12078
rect 12796 12014 12798 12066
rect 12850 12014 12852 12066
rect 12796 10834 12852 12014
rect 13580 11956 13636 11966
rect 12908 11508 12964 11518
rect 12908 11414 12964 11452
rect 13580 11394 13636 11900
rect 13580 11342 13582 11394
rect 13634 11342 13636 11394
rect 13580 11330 13636 11342
rect 13468 11284 13524 11294
rect 12796 10782 12798 10834
rect 12850 10782 12852 10834
rect 12796 10770 12852 10782
rect 13132 11282 13524 11284
rect 13132 11230 13470 11282
rect 13522 11230 13524 11282
rect 13132 11228 13524 11230
rect 13132 10722 13188 11228
rect 13468 11218 13524 11228
rect 13132 10670 13134 10722
rect 13186 10670 13188 10722
rect 13132 10658 13188 10670
rect 13692 10610 13748 12124
rect 13916 12114 13972 12124
rect 14364 11508 14420 12798
rect 14700 12290 14756 13020
rect 14700 12238 14702 12290
rect 14754 12238 14756 12290
rect 14700 12226 14756 12238
rect 13692 10558 13694 10610
rect 13746 10558 13748 10610
rect 11116 9986 11172 9996
rect 11340 9940 11396 9950
rect 11452 9940 11508 10444
rect 12460 10500 12516 10510
rect 12460 10406 12516 10444
rect 11340 9938 11508 9940
rect 11340 9886 11342 9938
rect 11394 9886 11508 9938
rect 11340 9884 11508 9886
rect 12572 9940 12628 9950
rect 11340 9874 11396 9884
rect 12572 9846 12628 9884
rect 13020 9940 13076 9950
rect 13020 9846 13076 9884
rect 13692 9940 13748 10558
rect 13692 9846 13748 9884
rect 13916 11394 13972 11406
rect 13916 11342 13918 11394
rect 13970 11342 13972 11394
rect 13916 11284 13972 11342
rect 13916 9938 13972 11228
rect 13916 9886 13918 9938
rect 13970 9886 13972 9938
rect 13916 9874 13972 9886
rect 14364 9716 14420 11452
rect 14924 11394 14980 14476
rect 15484 14530 15540 15092
rect 15484 14478 15486 14530
rect 15538 14478 15540 14530
rect 15484 14466 15540 14478
rect 15932 13972 15988 13982
rect 15932 13746 15988 13916
rect 16828 13972 16884 13982
rect 16828 13878 16884 13916
rect 16380 13860 16436 13870
rect 16380 13766 16436 13804
rect 17836 13860 17892 15092
rect 17948 15090 18004 15102
rect 18396 15092 18676 15148
rect 18732 15138 18788 15148
rect 19180 15314 19236 15372
rect 19180 15262 19182 15314
rect 19234 15262 19236 15314
rect 19180 15148 19236 15262
rect 19404 15314 19460 16156
rect 19404 15262 19406 15314
rect 19458 15262 19460 15314
rect 19404 15250 19460 15262
rect 19516 15316 19572 16380
rect 19628 15986 19684 16716
rect 19852 16706 19908 16716
rect 19628 15934 19630 15986
rect 19682 15934 19684 15986
rect 19628 15922 19684 15934
rect 19964 15876 20020 16828
rect 20188 16882 20244 16894
rect 20188 16830 20190 16882
rect 20242 16830 20244 16882
rect 20188 16100 20244 16830
rect 20244 16044 20356 16100
rect 20188 16034 20244 16044
rect 19964 15820 20244 15876
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20076 15540 20132 15550
rect 20188 15540 20244 15820
rect 20076 15538 20244 15540
rect 20076 15486 20078 15538
rect 20130 15486 20244 15538
rect 20076 15484 20244 15486
rect 20076 15474 20132 15484
rect 19628 15316 19684 15326
rect 20300 15316 20356 16044
rect 19516 15260 19628 15316
rect 19628 15222 19684 15260
rect 19852 15260 20356 15316
rect 19740 15204 19796 15214
rect 17948 15038 17950 15090
rect 18002 15038 18004 15090
rect 17948 14306 18004 15038
rect 17948 14254 17950 14306
rect 18002 14254 18004 14306
rect 17948 14242 18004 14254
rect 18508 14980 18564 14990
rect 17836 13766 17892 13804
rect 15932 13694 15934 13746
rect 15986 13694 15988 13746
rect 15932 13682 15988 13694
rect 18508 13300 18564 14924
rect 18620 14418 18676 15092
rect 19068 15092 19124 15102
rect 19180 15092 19572 15148
rect 19068 14868 19124 15036
rect 19068 14642 19124 14812
rect 19068 14590 19070 14642
rect 19122 14590 19124 14642
rect 19068 14578 19124 14590
rect 19292 14644 19348 14654
rect 18620 14366 18622 14418
rect 18674 14366 18676 14418
rect 18620 14084 18676 14366
rect 18620 14028 19124 14084
rect 19068 13746 19124 14028
rect 19068 13694 19070 13746
rect 19122 13694 19124 13746
rect 19068 13682 19124 13694
rect 19292 13970 19348 14588
rect 19292 13918 19294 13970
rect 19346 13918 19348 13970
rect 18844 13524 18900 13534
rect 18508 13244 18788 13300
rect 15260 13076 15316 13086
rect 15260 12982 15316 13020
rect 15596 13076 15652 13086
rect 14924 11342 14926 11394
rect 14978 11342 14980 11394
rect 14924 11330 14980 11342
rect 15596 11394 15652 13020
rect 18508 13076 18564 13114
rect 18508 13010 18564 13020
rect 18284 12850 18340 12862
rect 18284 12798 18286 12850
rect 18338 12798 18340 12850
rect 18284 12404 18340 12798
rect 18508 12852 18564 12862
rect 18508 12758 18564 12796
rect 17948 12402 18340 12404
rect 17948 12350 18286 12402
rect 18338 12350 18340 12402
rect 17948 12348 18340 12350
rect 16828 12124 17668 12180
rect 16828 12066 16884 12124
rect 16828 12014 16830 12066
rect 16882 12014 16884 12066
rect 16828 12002 16884 12014
rect 17388 11956 17444 11966
rect 17612 11956 17668 12124
rect 17948 12178 18004 12348
rect 18284 12338 18340 12348
rect 18732 12292 18788 13244
rect 18844 13186 18900 13468
rect 19292 13524 19348 13918
rect 19292 13458 19348 13468
rect 18844 13134 18846 13186
rect 18898 13134 18900 13186
rect 18844 13122 18900 13134
rect 19068 12964 19124 12974
rect 19404 12964 19460 12974
rect 19068 12962 19460 12964
rect 19068 12910 19070 12962
rect 19122 12910 19406 12962
rect 19458 12910 19460 12962
rect 19068 12908 19460 12910
rect 19516 12964 19572 15092
rect 19628 15092 19796 15148
rect 19628 14530 19684 15092
rect 19852 14754 19908 15260
rect 20412 15148 20468 17612
rect 20524 16100 20580 19966
rect 20860 19458 20916 20636
rect 21420 20580 21476 20590
rect 20972 20578 21476 20580
rect 20972 20526 21422 20578
rect 21474 20526 21476 20578
rect 20972 20524 21476 20526
rect 20972 20018 21028 20524
rect 21420 20514 21476 20524
rect 20972 19966 20974 20018
rect 21026 19966 21028 20018
rect 20972 19954 21028 19966
rect 20860 19406 20862 19458
rect 20914 19406 20916 19458
rect 20860 19394 20916 19406
rect 21420 19124 21476 19134
rect 21308 19012 21364 19022
rect 21308 18918 21364 18956
rect 21420 18788 21476 19068
rect 21196 18732 21476 18788
rect 21196 18004 21252 18732
rect 21420 18340 21476 18350
rect 21420 18246 21476 18284
rect 20748 17780 20804 17790
rect 20748 17444 20804 17724
rect 20748 16210 20804 17388
rect 20748 16158 20750 16210
rect 20802 16158 20804 16210
rect 20748 16146 20804 16158
rect 21084 16994 21140 17006
rect 21084 16942 21086 16994
rect 21138 16942 21140 16994
rect 21084 16212 21140 16942
rect 20524 16034 20580 16044
rect 19852 14702 19854 14754
rect 19906 14702 19908 14754
rect 19852 14690 19908 14702
rect 20300 15092 20468 15148
rect 20860 15426 20916 15438
rect 20860 15374 20862 15426
rect 20914 15374 20916 15426
rect 20860 15316 20916 15374
rect 21084 15316 21140 16156
rect 21196 15876 21252 17948
rect 21308 17892 21364 17902
rect 21308 17666 21364 17836
rect 21308 17614 21310 17666
rect 21362 17614 21364 17666
rect 21308 17602 21364 17614
rect 21532 17556 21588 21980
rect 22204 22148 22260 22158
rect 22204 21028 22260 22092
rect 22428 21700 22484 22206
rect 22428 21634 22484 21644
rect 22204 20962 22260 20972
rect 22316 21476 22372 21486
rect 22540 21476 22596 25228
rect 22652 25060 22708 26852
rect 22988 26740 23044 26750
rect 22652 24994 22708 25004
rect 22764 26290 22820 26302
rect 22764 26238 22766 26290
rect 22818 26238 22820 26290
rect 22652 24836 22708 24846
rect 22764 24836 22820 26238
rect 22988 26290 23044 26684
rect 23100 26514 23156 28028
rect 23100 26462 23102 26514
rect 23154 26462 23156 26514
rect 23100 26450 23156 26462
rect 23212 26404 23268 26414
rect 23212 26310 23268 26348
rect 22988 26238 22990 26290
rect 23042 26238 23044 26290
rect 22988 25732 23044 26238
rect 22876 25508 22932 25518
rect 22876 25414 22932 25452
rect 22988 25284 23044 25676
rect 23324 25620 23380 30156
rect 25228 30156 25620 30212
rect 25900 31554 25956 31566
rect 25900 31502 25902 31554
rect 25954 31502 25956 31554
rect 25900 30212 25956 31502
rect 26124 31220 26180 31230
rect 26124 31126 26180 31164
rect 26012 30996 26068 31006
rect 26012 30436 26068 30940
rect 26124 30436 26180 30446
rect 26012 30434 26180 30436
rect 26012 30382 26126 30434
rect 26178 30382 26180 30434
rect 26012 30380 26180 30382
rect 26124 30370 26180 30380
rect 24220 30098 24276 30110
rect 24556 30100 24612 30110
rect 24220 30046 24222 30098
rect 24274 30046 24276 30098
rect 24220 29988 24276 30046
rect 24220 29764 24276 29932
rect 24220 29698 24276 29708
rect 24444 30044 24556 30100
rect 24332 29540 24388 29550
rect 23660 29538 24388 29540
rect 23660 29486 24334 29538
rect 24386 29486 24388 29538
rect 23660 29484 24388 29486
rect 23660 28642 23716 29484
rect 24332 29474 24388 29484
rect 23660 28590 23662 28642
rect 23714 28590 23716 28642
rect 23660 28578 23716 28590
rect 23772 28084 23828 28094
rect 24332 28084 24388 28094
rect 24444 28084 24500 30044
rect 24556 30034 24612 30044
rect 25004 30100 25060 30110
rect 25004 30006 25060 30044
rect 24668 29988 24724 29998
rect 24668 29538 24724 29932
rect 25228 29540 25284 30156
rect 25900 30146 25956 30156
rect 25452 29988 25508 29998
rect 25788 29988 25844 29998
rect 25452 29986 25620 29988
rect 25452 29934 25454 29986
rect 25506 29934 25620 29986
rect 25452 29932 25620 29934
rect 25452 29922 25508 29932
rect 24668 29486 24670 29538
rect 24722 29486 24724 29538
rect 24668 29474 24724 29486
rect 25116 29484 25284 29540
rect 23660 28028 23772 28084
rect 23548 27970 23604 27982
rect 23548 27918 23550 27970
rect 23602 27918 23604 27970
rect 23436 27860 23492 27870
rect 23548 27860 23604 27918
rect 23436 27858 23604 27860
rect 23436 27806 23438 27858
rect 23490 27806 23604 27858
rect 23436 27804 23604 27806
rect 23436 27794 23492 27804
rect 23436 26292 23492 26302
rect 23436 26198 23492 26236
rect 22652 24834 22820 24836
rect 22652 24782 22654 24834
rect 22706 24782 22820 24834
rect 22652 24780 22820 24782
rect 22876 25228 23044 25284
rect 23100 25564 23380 25620
rect 22652 24770 22708 24780
rect 22876 24724 22932 25228
rect 22988 24836 23044 24846
rect 22988 24742 23044 24780
rect 22764 24668 22932 24724
rect 22652 23828 22708 23838
rect 22652 23154 22708 23772
rect 22652 23102 22654 23154
rect 22706 23102 22708 23154
rect 22652 23090 22708 23102
rect 22316 21474 22596 21476
rect 22316 21422 22318 21474
rect 22370 21422 22596 21474
rect 22316 21420 22596 21422
rect 21756 20692 21812 20702
rect 21756 20598 21812 20636
rect 22092 20690 22148 20702
rect 22092 20638 22094 20690
rect 22146 20638 22148 20690
rect 22092 20580 22148 20638
rect 22092 20514 22148 20524
rect 22204 19348 22260 19358
rect 22204 19254 22260 19292
rect 21644 18452 21700 18462
rect 21644 18358 21700 18396
rect 21756 18338 21812 18350
rect 21756 18286 21758 18338
rect 21810 18286 21812 18338
rect 21532 17332 21588 17500
rect 21532 17266 21588 17276
rect 21644 18116 21700 18126
rect 21308 16100 21364 16110
rect 21308 16006 21364 16044
rect 21196 15810 21252 15820
rect 21644 15540 21700 18060
rect 21756 16660 21812 18286
rect 21980 18340 22036 18350
rect 21980 18246 22036 18284
rect 21868 17778 21924 17790
rect 21868 17726 21870 17778
rect 21922 17726 21924 17778
rect 21868 17668 21924 17726
rect 21868 17602 21924 17612
rect 21980 16884 22036 16894
rect 22316 16884 22372 21420
rect 22652 20804 22708 20814
rect 22652 20710 22708 20748
rect 22764 19908 22820 24668
rect 22988 23826 23044 23838
rect 22988 23774 22990 23826
rect 23042 23774 23044 23826
rect 22876 23380 22932 23390
rect 22876 22820 22932 23324
rect 22988 23378 23044 23774
rect 22988 23326 22990 23378
rect 23042 23326 23044 23378
rect 22988 23314 23044 23326
rect 22876 22754 22932 22764
rect 23100 22708 23156 25564
rect 23660 25508 23716 28028
rect 23772 27990 23828 28028
rect 23884 28082 24500 28084
rect 23884 28030 24334 28082
rect 24386 28030 24500 28082
rect 23884 28028 24500 28030
rect 23884 27970 23940 28028
rect 24332 28018 24388 28028
rect 23884 27918 23886 27970
rect 23938 27918 23940 27970
rect 23884 27906 23940 27918
rect 24108 26852 24164 26862
rect 23884 26850 24164 26852
rect 23884 26798 24110 26850
rect 24162 26798 24164 26850
rect 23884 26796 24164 26798
rect 23884 26514 23940 26796
rect 24108 26786 24164 26796
rect 23884 26462 23886 26514
rect 23938 26462 23940 26514
rect 23884 26450 23940 26462
rect 23884 26292 23940 26302
rect 23772 26180 23828 26190
rect 23772 26086 23828 26124
rect 23772 25620 23828 25630
rect 23884 25620 23940 26236
rect 23996 26180 24052 26190
rect 24332 26180 24388 26190
rect 24052 26178 24388 26180
rect 24052 26126 24334 26178
rect 24386 26126 24388 26178
rect 24052 26124 24388 26126
rect 23996 26114 24052 26124
rect 24332 26114 24388 26124
rect 23828 25564 23940 25620
rect 24220 25732 24276 25742
rect 24220 25618 24276 25676
rect 24220 25566 24222 25618
rect 24274 25566 24276 25618
rect 23772 25526 23828 25564
rect 24220 25554 24276 25566
rect 23324 25394 23380 25406
rect 23324 25342 23326 25394
rect 23378 25342 23380 25394
rect 23324 25172 23380 25342
rect 23324 25106 23380 25116
rect 23660 24836 23716 25452
rect 24444 25396 24500 28028
rect 25116 28084 25172 29484
rect 25564 29428 25620 29932
rect 25788 29894 25844 29932
rect 24780 27860 24836 27870
rect 24780 27188 24836 27804
rect 24780 25506 24836 27132
rect 25004 27076 25060 27086
rect 25116 27076 25172 28028
rect 25004 27074 25172 27076
rect 25004 27022 25006 27074
rect 25058 27022 25172 27074
rect 25004 27020 25172 27022
rect 25228 29316 25284 29326
rect 25004 27010 25060 27020
rect 25228 26908 25284 29260
rect 25340 29204 25396 29214
rect 25340 29110 25396 29148
rect 25340 27748 25396 27758
rect 25340 27654 25396 27692
rect 25452 27188 25508 27198
rect 25452 27094 25508 27132
rect 25228 26852 25396 26908
rect 24780 25454 24782 25506
rect 24834 25454 24836 25506
rect 24780 25442 24836 25454
rect 25228 25508 25284 25518
rect 25228 25414 25284 25452
rect 24444 25330 24500 25340
rect 24444 25172 24500 25182
rect 24444 24946 24500 25116
rect 24444 24894 24446 24946
rect 24498 24894 24500 24946
rect 24444 24882 24500 24894
rect 23772 24836 23828 24846
rect 23660 24834 23828 24836
rect 23660 24782 23774 24834
rect 23826 24782 23828 24834
rect 23660 24780 23828 24782
rect 23324 24724 23380 24734
rect 23324 24722 23492 24724
rect 23324 24670 23326 24722
rect 23378 24670 23492 24722
rect 23324 24668 23492 24670
rect 23324 24658 23380 24668
rect 23212 24610 23268 24622
rect 23212 24558 23214 24610
rect 23266 24558 23268 24610
rect 23212 23940 23268 24558
rect 23436 24612 23492 24668
rect 23660 24612 23716 24622
rect 23436 24610 23716 24612
rect 23436 24558 23662 24610
rect 23714 24558 23716 24610
rect 23436 24556 23716 24558
rect 23660 24546 23716 24556
rect 23772 24612 23828 24780
rect 23996 24724 24052 24734
rect 23996 24630 24052 24668
rect 24332 24722 24388 24734
rect 24332 24670 24334 24722
rect 24386 24670 24388 24722
rect 23772 24546 23828 24556
rect 23212 23874 23268 23884
rect 23996 23940 24052 23950
rect 23996 23846 24052 23884
rect 24332 23828 24388 24670
rect 25228 24724 25284 24734
rect 25004 24612 25060 24622
rect 24332 23762 24388 23772
rect 24444 24498 24500 24510
rect 24444 24446 24446 24498
rect 24498 24446 24500 24498
rect 22988 22652 23156 22708
rect 23324 23714 23380 23726
rect 23324 23662 23326 23714
rect 23378 23662 23380 23714
rect 22876 20916 22932 20926
rect 22876 20822 22932 20860
rect 22988 20356 23044 22652
rect 23100 22484 23156 22494
rect 23100 22390 23156 22428
rect 23324 22370 23380 23662
rect 24220 23154 24276 23166
rect 24220 23102 24222 23154
rect 24274 23102 24276 23154
rect 24220 23044 24276 23102
rect 24220 22978 24276 22988
rect 23324 22318 23326 22370
rect 23378 22318 23380 22370
rect 23324 22306 23380 22318
rect 24444 22372 24500 24446
rect 25004 23938 25060 24556
rect 25004 23886 25006 23938
rect 25058 23886 25060 23938
rect 25004 23874 25060 23886
rect 25228 23266 25284 24668
rect 25228 23214 25230 23266
rect 25282 23214 25284 23266
rect 25228 23202 25284 23214
rect 24556 23156 24612 23166
rect 24556 23062 24612 23100
rect 24444 22306 24500 22316
rect 24668 23042 24724 23054
rect 24668 22990 24670 23042
rect 24722 22990 24724 23042
rect 23660 21700 23716 21710
rect 23548 21252 23604 21262
rect 23324 21028 23380 21038
rect 23100 20802 23156 20814
rect 23100 20750 23102 20802
rect 23154 20750 23156 20802
rect 23100 20468 23156 20750
rect 23324 20802 23380 20972
rect 23324 20750 23326 20802
rect 23378 20750 23380 20802
rect 23324 20738 23380 20750
rect 23548 20468 23604 21196
rect 23660 20580 23716 21644
rect 24220 21698 24276 21710
rect 24220 21646 24222 21698
rect 24274 21646 24276 21698
rect 24220 21588 24276 21646
rect 23884 21532 24276 21588
rect 24332 21586 24388 21598
rect 24332 21534 24334 21586
rect 24386 21534 24388 21586
rect 23660 20486 23716 20524
rect 23772 20692 23828 20702
rect 23100 20412 23604 20468
rect 23548 20356 23604 20412
rect 23548 20300 23716 20356
rect 22988 20290 23044 20300
rect 22764 19842 22820 19852
rect 23436 20242 23492 20254
rect 23436 20190 23438 20242
rect 23490 20190 23492 20242
rect 23100 19234 23156 19246
rect 23100 19182 23102 19234
rect 23154 19182 23156 19234
rect 22876 18564 22932 18574
rect 23100 18564 23156 19182
rect 23436 19124 23492 20190
rect 23436 19068 23604 19124
rect 22876 18562 23156 18564
rect 22876 18510 22878 18562
rect 22930 18510 23156 18562
rect 22876 18508 23156 18510
rect 22428 18338 22484 18350
rect 22428 18286 22430 18338
rect 22482 18286 22484 18338
rect 22428 18004 22484 18286
rect 22428 17938 22484 17948
rect 22764 17668 22820 17678
rect 22876 17668 22932 18508
rect 23212 18452 23268 18462
rect 23212 18450 23492 18452
rect 23212 18398 23214 18450
rect 23266 18398 23492 18450
rect 23212 18396 23492 18398
rect 23212 18386 23268 18396
rect 22820 17612 22932 17668
rect 22988 18340 23044 18350
rect 22764 17574 22820 17612
rect 22988 17108 23044 18284
rect 23212 18004 23268 18014
rect 23212 17778 23268 17948
rect 23212 17726 23214 17778
rect 23266 17726 23268 17778
rect 23212 17714 23268 17726
rect 22428 16884 22484 16894
rect 22316 16828 22428 16884
rect 21980 16790 22036 16828
rect 21756 16604 22036 16660
rect 21868 16098 21924 16110
rect 21868 16046 21870 16098
rect 21922 16046 21924 16098
rect 21756 15540 21812 15550
rect 21644 15538 21812 15540
rect 21644 15486 21758 15538
rect 21810 15486 21812 15538
rect 21644 15484 21812 15486
rect 21756 15474 21812 15484
rect 21756 15316 21812 15326
rect 21084 15314 21812 15316
rect 21084 15262 21758 15314
rect 21810 15262 21812 15314
rect 21084 15260 21812 15262
rect 20860 15148 20916 15260
rect 20860 15092 21252 15148
rect 19628 14478 19630 14530
rect 19682 14478 19684 14530
rect 19628 13858 19684 14478
rect 20188 14532 20244 14542
rect 20188 14438 20244 14476
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13806 19630 13858
rect 19682 13806 19684 13858
rect 19628 13794 19684 13806
rect 19740 12964 19796 12974
rect 19516 12962 19796 12964
rect 19516 12910 19742 12962
rect 19794 12910 19796 12962
rect 19516 12908 19796 12910
rect 19068 12898 19124 12908
rect 19404 12898 19460 12908
rect 19740 12898 19796 12908
rect 19628 12740 19684 12750
rect 20300 12740 20356 15092
rect 20524 14028 21140 14084
rect 20412 13748 20468 13758
rect 20524 13748 20580 14028
rect 21084 13970 21140 14028
rect 21084 13918 21086 13970
rect 21138 13918 21140 13970
rect 21084 13906 21140 13918
rect 20636 13860 20692 13870
rect 20636 13858 21028 13860
rect 20636 13806 20638 13858
rect 20690 13806 21028 13858
rect 20636 13804 21028 13806
rect 20636 13794 20692 13804
rect 20412 13746 20580 13748
rect 20412 13694 20414 13746
rect 20466 13694 20580 13746
rect 20412 13692 20580 13694
rect 20412 13682 20468 13692
rect 20412 13076 20468 13114
rect 20412 13010 20468 13020
rect 20524 12964 20580 12974
rect 19628 12738 20356 12740
rect 19628 12686 19630 12738
rect 19682 12686 20356 12738
rect 19628 12684 20356 12686
rect 18844 12292 18900 12302
rect 19292 12292 19348 12302
rect 18732 12290 19348 12292
rect 18732 12238 18846 12290
rect 18898 12238 19294 12290
rect 19346 12238 19348 12290
rect 18732 12236 19348 12238
rect 18844 12226 18900 12236
rect 17948 12126 17950 12178
rect 18002 12126 18004 12178
rect 17948 12114 18004 12126
rect 18396 12068 18452 12078
rect 18396 12066 18564 12068
rect 18396 12014 18398 12066
rect 18450 12014 18564 12066
rect 18396 12012 18564 12014
rect 18396 12002 18452 12012
rect 17724 11956 17780 11966
rect 17388 11954 17556 11956
rect 17388 11902 17390 11954
rect 17442 11902 17556 11954
rect 17388 11900 17556 11902
rect 17612 11954 17780 11956
rect 17612 11902 17726 11954
rect 17778 11902 17780 11954
rect 17612 11900 17780 11902
rect 17388 11890 17444 11900
rect 15596 11342 15598 11394
rect 15650 11342 15652 11394
rect 15596 11330 15652 11342
rect 16716 11732 16772 11742
rect 16716 10834 16772 11676
rect 16716 10782 16718 10834
rect 16770 10782 16772 10834
rect 16716 10770 16772 10782
rect 17500 10722 17556 11900
rect 17500 10670 17502 10722
rect 17554 10670 17556 10722
rect 17500 10658 17556 10670
rect 14476 10500 14532 10510
rect 14476 10498 14868 10500
rect 14476 10446 14478 10498
rect 14530 10446 14868 10498
rect 14476 10444 14868 10446
rect 14476 10434 14532 10444
rect 14812 10050 14868 10444
rect 14812 9998 14814 10050
rect 14866 9998 14868 10050
rect 14812 9986 14868 9998
rect 15372 9940 15428 9950
rect 15372 9846 15428 9884
rect 14476 9716 14532 9726
rect 14364 9714 14532 9716
rect 14364 9662 14478 9714
rect 14530 9662 14532 9714
rect 14364 9660 14532 9662
rect 14476 9650 14532 9660
rect 14028 9604 14084 9614
rect 14028 9602 14420 9604
rect 14028 9550 14030 9602
rect 14082 9550 14420 9602
rect 14028 9548 14420 9550
rect 14028 9538 14084 9548
rect 14364 9492 14420 9548
rect 14700 9602 14756 9614
rect 14700 9550 14702 9602
rect 14754 9550 14756 9602
rect 14700 9492 14756 9550
rect 14364 9436 14756 9492
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 17500 4340 17556 4350
rect 17724 4340 17780 11900
rect 18060 11508 18116 11518
rect 18060 11170 18116 11452
rect 18060 11118 18062 11170
rect 18114 11118 18116 11170
rect 18060 11106 18116 11118
rect 18508 11172 18564 12012
rect 18732 11954 18788 11966
rect 18732 11902 18734 11954
rect 18786 11902 18788 11954
rect 18732 11508 18788 11902
rect 18732 11442 18788 11452
rect 18620 11172 18676 11182
rect 19068 11172 19124 11182
rect 18508 11170 18676 11172
rect 18508 11118 18622 11170
rect 18674 11118 18676 11170
rect 18508 11116 18676 11118
rect 17836 10722 17892 10734
rect 17836 10670 17838 10722
rect 17890 10670 17892 10722
rect 17836 10612 17892 10670
rect 18172 10612 18228 10622
rect 17836 10610 18228 10612
rect 17836 10558 18174 10610
rect 18226 10558 18228 10610
rect 17836 10556 18228 10558
rect 18172 9042 18228 10556
rect 18172 8990 18174 9042
rect 18226 8990 18228 9042
rect 18172 7474 18228 8990
rect 18172 7422 18174 7474
rect 18226 7422 18228 7474
rect 18172 7410 18228 7422
rect 17500 4338 17780 4340
rect 17500 4286 17502 4338
rect 17554 4286 17780 4338
rect 17500 4284 17780 4286
rect 17500 4274 17556 4284
rect 17836 4226 17892 4238
rect 17836 4174 17838 4226
rect 17890 4174 17892 4226
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17836 3388 17892 4174
rect 17612 3332 17892 3388
rect 18172 3668 18228 3678
rect 16828 924 17108 980
rect 16828 800 16884 924
rect 17052 868 17108 924
rect 17052 812 17220 868
rect 16800 0 16912 800
rect 17164 756 17220 812
rect 17612 756 17668 3332
rect 18172 800 18228 3612
rect 18396 3444 18452 3454
rect 18508 3444 18564 11116
rect 18620 11106 18676 11116
rect 18732 11170 19124 11172
rect 18732 11118 19070 11170
rect 19122 11118 19124 11170
rect 18732 11116 19124 11118
rect 18732 10610 18788 11116
rect 19068 11106 19124 11116
rect 18732 10558 18734 10610
rect 18786 10558 18788 10610
rect 18732 10546 18788 10558
rect 18844 9940 18900 9950
rect 18844 9042 18900 9884
rect 19292 9940 19348 12236
rect 19628 11732 19684 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 20300 12292 20356 12684
rect 20300 12226 20356 12236
rect 20412 12850 20468 12862
rect 20412 12798 20414 12850
rect 20466 12798 20468 12850
rect 19964 12178 20020 12190
rect 19964 12126 19966 12178
rect 20018 12126 20020 12178
rect 19852 11954 19908 11966
rect 19852 11902 19854 11954
rect 19906 11902 19908 11954
rect 19852 11844 19908 11902
rect 19964 11956 20020 12126
rect 19964 11890 20020 11900
rect 19852 11778 19908 11788
rect 20412 11844 20468 12798
rect 19628 11666 19684 11676
rect 20412 11394 20468 11788
rect 20412 11342 20414 11394
rect 20466 11342 20468 11394
rect 20412 11330 20468 11342
rect 20524 11506 20580 12908
rect 20636 12964 20692 12974
rect 20636 12962 20804 12964
rect 20636 12910 20638 12962
rect 20690 12910 20804 12962
rect 20636 12908 20804 12910
rect 20636 12898 20692 12908
rect 20748 12404 20804 12908
rect 20972 12628 21028 13804
rect 21196 13746 21252 15092
rect 21196 13694 21198 13746
rect 21250 13694 21252 13746
rect 21196 13682 21252 13694
rect 21308 14980 21364 14990
rect 21308 14418 21364 14924
rect 21308 14366 21310 14418
rect 21362 14366 21364 14418
rect 21308 13860 21364 14366
rect 21532 14756 21588 14766
rect 21532 14306 21588 14700
rect 21532 14254 21534 14306
rect 21586 14254 21588 14306
rect 21532 14242 21588 14254
rect 21644 14420 21700 14430
rect 21084 13522 21140 13534
rect 21084 13470 21086 13522
rect 21138 13470 21140 13522
rect 21084 12964 21140 13470
rect 21308 13076 21364 13804
rect 21644 13746 21700 14364
rect 21644 13694 21646 13746
rect 21698 13694 21700 13746
rect 21644 13682 21700 13694
rect 21420 13636 21476 13646
rect 21756 13636 21812 15260
rect 21868 14756 21924 16046
rect 21868 14690 21924 14700
rect 21868 14532 21924 14542
rect 21980 14532 22036 16604
rect 22092 15316 22148 15326
rect 22092 15222 22148 15260
rect 21868 14530 22036 14532
rect 21868 14478 21870 14530
rect 21922 14478 22036 14530
rect 21868 14476 22036 14478
rect 22204 14532 22260 14542
rect 21868 14466 21924 14476
rect 22204 14438 22260 14476
rect 22428 13972 22484 16828
rect 22988 15148 23044 17052
rect 23100 17332 23156 17342
rect 23100 16994 23156 17276
rect 23100 16942 23102 16994
rect 23154 16942 23156 16994
rect 23100 16930 23156 16942
rect 23324 15316 23380 15326
rect 23324 15222 23380 15260
rect 22764 15092 23044 15148
rect 23212 15202 23268 15214
rect 23212 15150 23214 15202
rect 23266 15150 23268 15202
rect 22540 14644 22596 14654
rect 22540 14418 22596 14588
rect 22540 14366 22542 14418
rect 22594 14366 22596 14418
rect 22540 14354 22596 14366
rect 21980 13916 22372 13972
rect 21756 13580 21924 13636
rect 21420 13542 21476 13580
rect 21644 13076 21700 13086
rect 21308 13074 21700 13076
rect 21308 13022 21646 13074
rect 21698 13022 21700 13074
rect 21308 13020 21700 13022
rect 21644 13010 21700 13020
rect 21084 12898 21140 12908
rect 21868 12852 21924 13580
rect 21868 12786 21924 12796
rect 20972 12572 21140 12628
rect 20972 12404 21028 12414
rect 20748 12402 21028 12404
rect 20748 12350 20974 12402
rect 21026 12350 21028 12402
rect 20748 12348 21028 12350
rect 20860 12180 20916 12190
rect 20860 12086 20916 12124
rect 20524 11454 20526 11506
rect 20578 11454 20580 11506
rect 19404 11284 19460 11294
rect 19740 11284 19796 11294
rect 19404 11282 19796 11284
rect 19404 11230 19406 11282
rect 19458 11230 19742 11282
rect 19794 11230 19796 11282
rect 19404 11228 19796 11230
rect 19404 11218 19460 11228
rect 19740 11218 19796 11228
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19740 10052 19796 10062
rect 19740 9958 19796 9996
rect 19628 9940 19684 9950
rect 19292 9938 19684 9940
rect 19292 9886 19294 9938
rect 19346 9886 19630 9938
rect 19682 9886 19684 9938
rect 19292 9884 19684 9886
rect 19292 9874 19348 9884
rect 19628 9604 19684 9884
rect 20524 9938 20580 11454
rect 20524 9886 20526 9938
rect 20578 9886 20580 9938
rect 20524 9874 20580 9886
rect 20748 12066 20804 12078
rect 20748 12014 20750 12066
rect 20802 12014 20804 12066
rect 20748 9828 20804 12014
rect 20972 11284 21028 12348
rect 20972 11218 21028 11228
rect 20972 10722 21028 10734
rect 20972 10670 20974 10722
rect 21026 10670 21028 10722
rect 20972 10052 21028 10670
rect 20972 9986 21028 9996
rect 20636 9772 20748 9828
rect 19628 9538 19684 9548
rect 20524 9716 20580 9726
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 18844 8990 18846 9042
rect 18898 8990 18900 9042
rect 18844 8978 18900 8990
rect 20412 8260 20468 8270
rect 20524 8260 20580 9660
rect 20636 8370 20692 9772
rect 20748 9734 20804 9772
rect 20636 8318 20638 8370
rect 20690 8318 20692 8370
rect 20636 8306 20692 8318
rect 20412 8258 20580 8260
rect 20412 8206 20414 8258
rect 20466 8206 20580 8258
rect 20412 8204 20580 8206
rect 20412 8194 20468 8204
rect 19404 8148 19460 8158
rect 19740 8148 19796 8158
rect 19404 8146 19796 8148
rect 19404 8094 19406 8146
rect 19458 8094 19742 8146
rect 19794 8094 19796 8146
rect 19404 8092 19796 8094
rect 19404 8082 19460 8092
rect 19740 8082 19796 8092
rect 19068 8036 19124 8046
rect 18844 8034 19124 8036
rect 18844 7982 19070 8034
rect 19122 7982 19124 8034
rect 18844 7980 19124 7982
rect 18844 7474 18900 7980
rect 19068 7970 19124 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 18844 7422 18846 7474
rect 18898 7422 18900 7474
rect 18844 7410 18900 7422
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 18844 3668 18900 3678
rect 18844 3574 18900 3612
rect 18396 3442 18564 3444
rect 18396 3390 18398 3442
rect 18450 3390 18564 3442
rect 18396 3388 18564 3390
rect 21084 3444 21140 12572
rect 21980 12292 22036 13916
rect 22204 13746 22260 13758
rect 22204 13694 22206 13746
rect 22258 13694 22260 13746
rect 22092 12964 22148 12974
rect 22092 12870 22148 12908
rect 21980 12290 22148 12292
rect 21980 12238 21982 12290
rect 22034 12238 22148 12290
rect 21980 12236 22148 12238
rect 21980 12226 22036 12236
rect 21868 11284 21924 11294
rect 21868 11190 21924 11228
rect 22092 10052 22148 12236
rect 22204 12180 22260 13694
rect 22316 13748 22372 13916
rect 22428 13906 22484 13916
rect 22652 13860 22708 13870
rect 22540 13858 22708 13860
rect 22540 13806 22654 13858
rect 22706 13806 22708 13858
rect 22540 13804 22708 13806
rect 22540 13748 22596 13804
rect 22652 13794 22708 13804
rect 22316 13692 22596 13748
rect 22652 12852 22708 12862
rect 22260 12124 22484 12180
rect 22204 12086 22260 12124
rect 22204 10500 22260 10510
rect 22204 10406 22260 10444
rect 21644 9996 22148 10052
rect 21644 9940 21700 9996
rect 22092 9940 22148 9996
rect 22316 9940 22372 9950
rect 22092 9938 22372 9940
rect 22092 9886 22318 9938
rect 22370 9886 22372 9938
rect 22092 9884 22372 9886
rect 21644 9846 21700 9884
rect 22316 9874 22372 9884
rect 21308 9828 21364 9838
rect 21308 9734 21364 9772
rect 21868 9828 21924 9838
rect 21420 9604 21476 9614
rect 21308 9266 21364 9278
rect 21308 9214 21310 9266
rect 21362 9214 21364 9266
rect 21308 8482 21364 9214
rect 21308 8430 21310 8482
rect 21362 8430 21364 8482
rect 21308 8418 21364 8430
rect 21420 8370 21476 9548
rect 21868 9268 21924 9772
rect 22428 9826 22484 12124
rect 22652 11506 22708 12796
rect 22764 12068 22820 15092
rect 22876 14418 22932 14430
rect 22876 14366 22878 14418
rect 22930 14366 22932 14418
rect 22876 13074 22932 14366
rect 23212 14420 23268 15150
rect 23436 15148 23492 18396
rect 23548 18450 23604 19068
rect 23660 18676 23716 20300
rect 23772 19458 23828 20636
rect 23884 19796 23940 21532
rect 24220 21364 24276 21374
rect 24220 21270 24276 21308
rect 24220 20916 24276 20926
rect 24108 20860 24220 20916
rect 23996 20804 24052 20814
rect 23996 20244 24052 20748
rect 23996 20178 24052 20188
rect 23996 19796 24052 19806
rect 23884 19794 24052 19796
rect 23884 19742 23998 19794
rect 24050 19742 24052 19794
rect 23884 19740 24052 19742
rect 23772 19406 23774 19458
rect 23826 19406 23828 19458
rect 23772 19394 23828 19406
rect 23996 19236 24052 19740
rect 24108 19684 24164 20860
rect 24220 20822 24276 20860
rect 24108 19618 24164 19628
rect 24220 20356 24276 20366
rect 24220 20130 24276 20300
rect 24220 20078 24222 20130
rect 24274 20078 24276 20130
rect 24108 19236 24164 19246
rect 23996 19180 24108 19236
rect 24220 19236 24276 20078
rect 24332 19460 24388 21534
rect 24668 21140 24724 22990
rect 24668 21074 24724 21084
rect 24780 23044 24836 23054
rect 24668 20916 24724 20926
rect 24780 20916 24836 22988
rect 25340 22036 25396 26852
rect 25452 25396 25508 25406
rect 25452 24948 25508 25340
rect 25564 25284 25620 29372
rect 26012 29764 26068 29774
rect 25788 29316 25844 29326
rect 25788 29222 25844 29260
rect 25900 29204 25956 29214
rect 25900 28530 25956 29148
rect 25900 28478 25902 28530
rect 25954 28478 25956 28530
rect 25900 28466 25956 28478
rect 25900 27076 25956 27086
rect 25900 26982 25956 27020
rect 25564 25218 25620 25228
rect 25900 24948 25956 24958
rect 25452 24946 25844 24948
rect 25452 24894 25454 24946
rect 25506 24894 25844 24946
rect 25452 24892 25844 24894
rect 25452 24882 25508 24892
rect 25788 24834 25844 24892
rect 25900 24854 25956 24892
rect 25788 24782 25790 24834
rect 25842 24782 25844 24834
rect 25788 24770 25844 24782
rect 25900 24724 25956 24734
rect 25900 23938 25956 24668
rect 25900 23886 25902 23938
rect 25954 23886 25956 23938
rect 25900 23874 25956 23886
rect 26012 23828 26068 29708
rect 26236 29652 26292 32396
rect 26348 31892 26404 31902
rect 26348 31798 26404 31836
rect 26572 31780 26628 31790
rect 26572 31686 26628 31724
rect 26684 30996 26740 35420
rect 27020 35252 27076 35756
rect 27132 35746 27188 35756
rect 27356 35698 27412 35868
rect 27356 35646 27358 35698
rect 27410 35646 27412 35698
rect 27356 35634 27412 35646
rect 27580 35308 27636 36316
rect 27692 36278 27748 36316
rect 27804 36036 27860 37212
rect 27916 37202 27972 37212
rect 28028 36484 28084 36494
rect 28252 36484 28308 36494
rect 28028 36482 28308 36484
rect 28028 36430 28030 36482
rect 28082 36430 28254 36482
rect 28306 36430 28308 36482
rect 28028 36428 28308 36430
rect 28028 36418 28084 36428
rect 28252 36418 28308 36428
rect 26796 35196 27076 35252
rect 27132 35252 27636 35308
rect 27692 35980 27860 36036
rect 28476 36372 28532 36382
rect 26796 34132 26852 35196
rect 27132 35140 27188 35252
rect 27020 35084 27188 35140
rect 26908 34802 26964 34814
rect 26908 34750 26910 34802
rect 26962 34750 26964 34802
rect 26908 34692 26964 34750
rect 27020 34692 27076 35084
rect 27132 34916 27188 34926
rect 27132 34914 27636 34916
rect 27132 34862 27134 34914
rect 27186 34862 27636 34914
rect 27132 34860 27636 34862
rect 27132 34850 27188 34860
rect 27244 34692 27300 34702
rect 27020 34690 27300 34692
rect 27020 34638 27246 34690
rect 27298 34638 27300 34690
rect 27020 34636 27300 34638
rect 26908 34626 26964 34636
rect 27244 34626 27300 34636
rect 27356 34692 27412 34702
rect 27356 34598 27412 34636
rect 27468 34690 27524 34702
rect 27468 34638 27470 34690
rect 27522 34638 27524 34690
rect 27244 34356 27300 34366
rect 27132 34132 27188 34142
rect 26796 34076 27132 34132
rect 27132 33908 27188 34076
rect 27132 33842 27188 33852
rect 27244 33684 27300 34300
rect 27356 34130 27412 34142
rect 27356 34078 27358 34130
rect 27410 34078 27412 34130
rect 27356 33796 27412 34078
rect 27356 33730 27412 33740
rect 26908 33628 27300 33684
rect 26908 33346 26964 33628
rect 27132 33460 27188 33470
rect 26908 33294 26910 33346
rect 26962 33294 26964 33346
rect 26908 33282 26964 33294
rect 27020 33458 27188 33460
rect 27020 33406 27134 33458
rect 27186 33406 27188 33458
rect 27020 33404 27188 33406
rect 26908 32676 26964 32686
rect 27020 32676 27076 33404
rect 27132 33394 27188 33404
rect 26964 32620 27076 32676
rect 27132 32786 27188 32798
rect 27132 32734 27134 32786
rect 27186 32734 27188 32786
rect 26908 32582 26964 32620
rect 27020 31892 27076 31902
rect 26796 31780 26852 31790
rect 26796 31554 26852 31724
rect 27020 31778 27076 31836
rect 27020 31726 27022 31778
rect 27074 31726 27076 31778
rect 26908 31668 26964 31678
rect 26908 31574 26964 31612
rect 26796 31502 26798 31554
rect 26850 31502 26852 31554
rect 26796 31220 26852 31502
rect 26796 31154 26852 31164
rect 26796 30996 26852 31006
rect 26740 30994 26852 30996
rect 26740 30942 26798 30994
rect 26850 30942 26852 30994
rect 26740 30940 26852 30942
rect 26348 30100 26404 30110
rect 26348 30006 26404 30044
rect 26572 30100 26628 30110
rect 26236 29596 26516 29652
rect 26348 29428 26404 29438
rect 26348 29334 26404 29372
rect 26348 28308 26404 28318
rect 26348 28082 26404 28252
rect 26348 28030 26350 28082
rect 26402 28030 26404 28082
rect 26236 27076 26292 27114
rect 26236 27010 26292 27020
rect 26348 26908 26404 28030
rect 26236 26852 26404 26908
rect 26460 26852 26516 29596
rect 26572 28644 26628 30044
rect 26684 28866 26740 30940
rect 26796 30930 26852 30940
rect 27020 30882 27076 31726
rect 27020 30830 27022 30882
rect 27074 30830 27076 30882
rect 27020 30818 27076 30830
rect 27132 30660 27188 32734
rect 27244 32562 27300 33628
rect 27468 33460 27524 34638
rect 27580 34242 27636 34860
rect 27580 34190 27582 34242
rect 27634 34190 27636 34242
rect 27580 34178 27636 34190
rect 27580 33460 27636 33470
rect 27468 33458 27636 33460
rect 27468 33406 27582 33458
rect 27634 33406 27636 33458
rect 27468 33404 27636 33406
rect 27580 33394 27636 33404
rect 27244 32510 27246 32562
rect 27298 32510 27300 32562
rect 27244 31556 27300 32510
rect 27356 33124 27412 33134
rect 27356 32562 27412 33068
rect 27356 32510 27358 32562
rect 27410 32510 27412 32562
rect 27356 32452 27412 32510
rect 27356 32386 27412 32396
rect 27692 32900 27748 35980
rect 28364 35924 28420 35934
rect 28364 35830 28420 35868
rect 28476 35700 28532 36316
rect 28588 36372 28644 36382
rect 28700 36372 28756 37324
rect 28588 36370 28756 36372
rect 28588 36318 28590 36370
rect 28642 36318 28756 36370
rect 28588 36316 28756 36318
rect 28588 36306 28644 36316
rect 28140 35644 28532 35700
rect 27916 35588 27972 35598
rect 27916 35494 27972 35532
rect 28140 34802 28196 35644
rect 28140 34750 28142 34802
rect 28194 34750 28196 34802
rect 28140 34738 28196 34750
rect 28252 34802 28308 34814
rect 28252 34750 28254 34802
rect 28306 34750 28308 34802
rect 27916 34692 27972 34702
rect 27804 34690 27972 34692
rect 27804 34638 27918 34690
rect 27970 34638 27972 34690
rect 27804 34636 27972 34638
rect 27804 33572 27860 34636
rect 27916 34626 27972 34636
rect 27916 34356 27972 34366
rect 28252 34356 28308 34750
rect 27916 34242 27972 34300
rect 27916 34190 27918 34242
rect 27970 34190 27972 34242
rect 27916 34178 27972 34190
rect 28028 34300 28308 34356
rect 28364 34692 28420 34702
rect 28028 34244 28084 34300
rect 28028 34130 28084 34188
rect 28028 34078 28030 34130
rect 28082 34078 28084 34130
rect 28028 34066 28084 34078
rect 28140 34132 28196 34142
rect 27804 33506 27860 33516
rect 27916 33796 27972 33806
rect 27916 33570 27972 33740
rect 27916 33518 27918 33570
rect 27970 33518 27972 33570
rect 27916 33506 27972 33518
rect 28140 33234 28196 34076
rect 28140 33182 28142 33234
rect 28194 33182 28196 33234
rect 28140 33170 28196 33182
rect 28252 33458 28308 33470
rect 28252 33406 28254 33458
rect 28306 33406 28308 33458
rect 27692 32844 28084 32900
rect 27692 31892 27748 32844
rect 27916 32676 27972 32686
rect 27692 31826 27748 31836
rect 27804 32674 27972 32676
rect 27804 32622 27918 32674
rect 27970 32622 27972 32674
rect 27804 32620 27972 32622
rect 27804 31780 27860 32620
rect 27916 32610 27972 32620
rect 28028 32676 28084 32844
rect 28028 32582 28084 32620
rect 28140 32452 28196 32462
rect 27804 31714 27860 31724
rect 27916 32338 27972 32350
rect 27916 32286 27918 32338
rect 27970 32286 27972 32338
rect 27916 31778 27972 32286
rect 28028 31892 28084 31902
rect 28028 31798 28084 31836
rect 27916 31726 27918 31778
rect 27970 31726 27972 31778
rect 27916 31714 27972 31726
rect 28140 31778 28196 32396
rect 28140 31726 28142 31778
rect 28194 31726 28196 31778
rect 28140 31714 28196 31726
rect 28252 31780 28308 33406
rect 27580 31668 27636 31678
rect 27580 31574 27636 31612
rect 27244 31490 27300 31500
rect 27468 30884 27524 30894
rect 27468 30790 27524 30828
rect 27804 30884 27860 30894
rect 27804 30882 28084 30884
rect 27804 30830 27806 30882
rect 27858 30830 28084 30882
rect 27804 30828 28084 30830
rect 27804 30818 27860 30828
rect 27132 30604 27524 30660
rect 27468 30210 27524 30604
rect 27468 30158 27470 30210
rect 27522 30158 27524 30210
rect 27468 30146 27524 30158
rect 27916 30212 27972 30222
rect 27916 30118 27972 30156
rect 26908 30100 26964 30110
rect 26908 30006 26964 30044
rect 27356 30098 27412 30110
rect 27356 30046 27358 30098
rect 27410 30046 27412 30098
rect 27356 29428 27412 30046
rect 27804 30100 27860 30110
rect 27356 29372 27636 29428
rect 26684 28814 26686 28866
rect 26738 28814 26740 28866
rect 26684 28802 26740 28814
rect 27356 28756 27412 28766
rect 27356 28662 27412 28700
rect 27580 28754 27636 29372
rect 27580 28702 27582 28754
rect 27634 28702 27636 28754
rect 27580 28690 27636 28702
rect 27804 28756 27860 30044
rect 27916 28756 27972 28766
rect 27804 28754 27972 28756
rect 27804 28702 27918 28754
rect 27970 28702 27972 28754
rect 27804 28700 27972 28702
rect 27916 28690 27972 28700
rect 26572 28588 26964 28644
rect 26572 27860 26628 27870
rect 26572 27766 26628 27804
rect 26684 27748 26740 27758
rect 26684 27412 26740 27692
rect 26908 27636 26964 28588
rect 27020 28532 27076 28542
rect 27020 28438 27076 28476
rect 27804 28532 27860 28542
rect 27804 28438 27860 28476
rect 28028 28530 28084 30828
rect 28252 30882 28308 31724
rect 28252 30830 28254 30882
rect 28306 30830 28308 30882
rect 28252 30818 28308 30830
rect 28028 28478 28030 28530
rect 28082 28478 28084 28530
rect 28028 28466 28084 28478
rect 27244 28028 27860 28084
rect 27244 27858 27300 28028
rect 27244 27806 27246 27858
rect 27298 27806 27300 27858
rect 27244 27794 27300 27806
rect 27580 27860 27636 27870
rect 26908 27580 27524 27636
rect 26684 27186 26740 27356
rect 26684 27134 26686 27186
rect 26738 27134 26740 27186
rect 26684 26908 26740 27134
rect 27468 27188 27524 27580
rect 27468 27094 27524 27132
rect 26684 26852 26852 26908
rect 26236 26516 26292 26852
rect 26460 26786 26516 26796
rect 26236 24948 26292 26460
rect 26348 26292 26404 26302
rect 26684 26292 26740 26302
rect 26348 26290 26740 26292
rect 26348 26238 26350 26290
rect 26402 26238 26686 26290
rect 26738 26238 26740 26290
rect 26348 26236 26740 26238
rect 26348 26226 26404 26236
rect 26684 26180 26740 26236
rect 26684 26114 26740 26124
rect 26796 25732 26852 26852
rect 27356 26292 27412 26302
rect 27356 26178 27412 26236
rect 27356 26126 27358 26178
rect 27410 26126 27412 26178
rect 27356 26114 27412 26126
rect 26684 25676 26852 25732
rect 26236 24892 26404 24948
rect 26124 24834 26180 24846
rect 26124 24782 26126 24834
rect 26178 24782 26180 24834
rect 26124 24724 26180 24782
rect 26236 24724 26292 24734
rect 26124 24722 26292 24724
rect 26124 24670 26238 24722
rect 26290 24670 26292 24722
rect 26124 24668 26292 24670
rect 26236 24658 26292 24668
rect 26012 23762 26068 23772
rect 24668 20914 24836 20916
rect 24668 20862 24670 20914
rect 24722 20862 24836 20914
rect 24668 20860 24836 20862
rect 25228 21980 25396 22036
rect 25452 23154 25508 23166
rect 25900 23156 25956 23166
rect 25452 23102 25454 23154
rect 25506 23102 25508 23154
rect 25452 22148 25508 23102
rect 25676 23154 25956 23156
rect 25676 23102 25902 23154
rect 25954 23102 25956 23154
rect 25676 23100 25956 23102
rect 25676 23044 25732 23100
rect 25900 23090 25956 23100
rect 25676 22482 25732 22988
rect 26236 23044 26292 23054
rect 25900 22932 25956 22942
rect 25900 22838 25956 22876
rect 25676 22430 25678 22482
rect 25730 22430 25732 22482
rect 25676 22418 25732 22430
rect 25788 22372 25844 22382
rect 25788 22278 25844 22316
rect 26236 22370 26292 22988
rect 26236 22318 26238 22370
rect 26290 22318 26292 22370
rect 26236 22306 26292 22318
rect 24668 20850 24724 20860
rect 24444 20580 24500 20590
rect 24444 20242 24500 20524
rect 25228 20468 25284 21980
rect 25340 21812 25396 21822
rect 25340 21718 25396 21756
rect 25452 21252 25508 22092
rect 25452 21186 25508 21196
rect 25676 21586 25732 21598
rect 25676 21534 25678 21586
rect 25730 21534 25732 21586
rect 25452 20914 25508 20926
rect 25452 20862 25454 20914
rect 25506 20862 25508 20914
rect 25228 20412 25396 20468
rect 24444 20190 24446 20242
rect 24498 20190 24500 20242
rect 24444 20178 24500 20190
rect 25228 20244 25284 20254
rect 25228 20150 25284 20188
rect 24780 20020 24836 20030
rect 24780 19926 24836 19964
rect 24556 19796 24612 19806
rect 24556 19702 24612 19740
rect 25340 19684 25396 20412
rect 25452 20132 25508 20862
rect 25452 20020 25508 20076
rect 25564 20020 25620 20030
rect 25452 20018 25620 20020
rect 25452 19966 25566 20018
rect 25618 19966 25620 20018
rect 25452 19964 25620 19966
rect 25564 19954 25620 19964
rect 25340 19628 25620 19684
rect 24332 19394 24388 19404
rect 24668 19572 24724 19582
rect 24220 19180 24612 19236
rect 24108 19142 24164 19180
rect 24220 18676 24276 18686
rect 23660 18674 24276 18676
rect 23660 18622 24222 18674
rect 24274 18622 24276 18674
rect 23660 18620 24276 18622
rect 24220 18610 24276 18620
rect 24556 18674 24612 19180
rect 24556 18622 24558 18674
rect 24610 18622 24612 18674
rect 23548 18398 23550 18450
rect 23602 18398 23604 18450
rect 23548 18386 23604 18398
rect 23660 18338 23716 18350
rect 23660 18286 23662 18338
rect 23714 18286 23716 18338
rect 23660 18004 23716 18286
rect 23660 17938 23716 17948
rect 23772 18228 23828 18238
rect 23884 18228 23940 18238
rect 23828 18226 23940 18228
rect 23828 18174 23886 18226
rect 23938 18174 23940 18226
rect 23828 18172 23940 18174
rect 23772 17106 23828 18172
rect 23884 18162 23940 18172
rect 24556 18116 24612 18622
rect 24668 19234 24724 19516
rect 25340 19460 25396 19470
rect 25340 19366 25396 19404
rect 24668 19182 24670 19234
rect 24722 19182 24724 19234
rect 24668 18226 24724 19182
rect 24892 19124 24948 19134
rect 24892 19030 24948 19068
rect 24668 18174 24670 18226
rect 24722 18174 24724 18226
rect 24668 18162 24724 18174
rect 25452 18450 25508 18462
rect 25452 18398 25454 18450
rect 25506 18398 25508 18450
rect 24556 18050 24612 18060
rect 24108 18004 24164 18014
rect 23772 17054 23774 17106
rect 23826 17054 23828 17106
rect 23772 17042 23828 17054
rect 23996 17666 24052 17678
rect 23996 17614 23998 17666
rect 24050 17614 24052 17666
rect 23996 16100 24052 17614
rect 24108 17106 24164 17948
rect 24108 17054 24110 17106
rect 24162 17054 24164 17106
rect 24108 17042 24164 17054
rect 24668 17666 24724 17678
rect 24668 17614 24670 17666
rect 24722 17614 24724 17666
rect 24556 16996 24612 17006
rect 24556 16902 24612 16940
rect 23996 16034 24052 16044
rect 24444 16658 24500 16670
rect 24444 16606 24446 16658
rect 24498 16606 24500 16658
rect 24444 15874 24500 16606
rect 24444 15822 24446 15874
rect 24498 15822 24500 15874
rect 24444 15810 24500 15822
rect 24668 15540 24724 17614
rect 25452 17668 25508 18398
rect 25564 18340 25620 19628
rect 25676 19458 25732 21534
rect 26012 21140 26068 21150
rect 25788 20802 25844 20814
rect 25788 20750 25790 20802
rect 25842 20750 25844 20802
rect 25788 20468 25844 20750
rect 25844 20412 25956 20468
rect 25788 20402 25844 20412
rect 25676 19406 25678 19458
rect 25730 19406 25732 19458
rect 25676 19394 25732 19406
rect 25788 19906 25844 19918
rect 25788 19854 25790 19906
rect 25842 19854 25844 19906
rect 25676 19236 25732 19246
rect 25676 19142 25732 19180
rect 25788 18452 25844 19854
rect 25900 19236 25956 20412
rect 26012 19236 26068 21084
rect 26236 20132 26292 20142
rect 26236 19908 26292 20076
rect 26236 19842 26292 19852
rect 26124 19794 26180 19806
rect 26124 19742 26126 19794
rect 26178 19742 26180 19794
rect 26124 19460 26180 19742
rect 26124 19394 26180 19404
rect 26124 19236 26180 19246
rect 26012 19234 26180 19236
rect 26012 19182 26126 19234
rect 26178 19182 26180 19234
rect 26012 19180 26180 19182
rect 25900 19170 25956 19180
rect 26124 19170 26180 19180
rect 26348 19234 26404 24892
rect 26684 24946 26740 25676
rect 26684 24894 26686 24946
rect 26738 24894 26740 24946
rect 26684 24724 26740 24894
rect 26796 25508 26852 25518
rect 26796 24946 26852 25452
rect 27468 25282 27524 25294
rect 27468 25230 27470 25282
rect 27522 25230 27524 25282
rect 26796 24894 26798 24946
rect 26850 24894 26852 24946
rect 26796 24882 26852 24894
rect 27356 24948 27412 24958
rect 27468 24948 27524 25230
rect 27356 24946 27524 24948
rect 27356 24894 27358 24946
rect 27410 24894 27524 24946
rect 27356 24892 27524 24894
rect 27356 24882 27412 24892
rect 27244 24836 27300 24846
rect 27244 24742 27300 24780
rect 26684 24658 26740 24668
rect 26908 24724 26964 24734
rect 26908 24722 27188 24724
rect 26908 24670 26910 24722
rect 26962 24670 27188 24722
rect 26908 24668 27188 24670
rect 26908 24658 26964 24668
rect 27132 24050 27188 24668
rect 27580 24722 27636 27804
rect 27804 26962 27860 28028
rect 27804 26910 27806 26962
rect 27858 26910 27860 26962
rect 27804 26898 27860 26910
rect 28140 26964 28196 27002
rect 28140 26898 28196 26908
rect 28364 26292 28420 34636
rect 28476 34130 28532 35644
rect 28476 34078 28478 34130
rect 28530 34078 28532 34130
rect 28476 34066 28532 34078
rect 28700 35028 28756 36316
rect 28924 35922 28980 37438
rect 29484 37380 29540 37772
rect 29708 37762 29764 37772
rect 29820 37826 29988 37828
rect 29820 37774 29934 37826
rect 29986 37774 29988 37826
rect 29820 37772 29988 37774
rect 29484 37314 29540 37324
rect 29596 37492 29652 37502
rect 29820 37492 29876 37772
rect 29932 37762 29988 37772
rect 31276 37826 31332 37838
rect 31276 37774 31278 37826
rect 31330 37774 31332 37826
rect 29596 37490 29876 37492
rect 29596 37438 29598 37490
rect 29650 37438 29876 37490
rect 29596 37436 29876 37438
rect 30268 37492 30324 37502
rect 29036 36932 29092 36942
rect 29036 36482 29092 36876
rect 29036 36430 29038 36482
rect 29090 36430 29092 36482
rect 29036 36418 29092 36430
rect 29596 36372 29652 37436
rect 29820 37268 29876 37278
rect 29820 37174 29876 37212
rect 30268 37266 30324 37436
rect 30268 37214 30270 37266
rect 30322 37214 30324 37266
rect 30268 37202 30324 37214
rect 31164 37266 31220 37278
rect 31164 37214 31166 37266
rect 31218 37214 31220 37266
rect 30828 37154 30884 37166
rect 30828 37102 30830 37154
rect 30882 37102 30884 37154
rect 29820 36932 29876 36942
rect 29708 36484 29764 36494
rect 29708 36390 29764 36428
rect 29596 36306 29652 36316
rect 28924 35870 28926 35922
rect 28978 35870 28980 35922
rect 28924 35858 28980 35870
rect 29372 36260 29428 36270
rect 29372 35922 29428 36204
rect 29372 35870 29374 35922
rect 29426 35870 29428 35922
rect 29372 35858 29428 35870
rect 29820 35922 29876 36876
rect 30828 36708 30884 37102
rect 30492 36652 30884 36708
rect 30940 37042 30996 37054
rect 30940 36990 30942 37042
rect 30994 36990 30996 37042
rect 30268 36260 30324 36270
rect 30324 36204 30436 36260
rect 30268 36194 30324 36204
rect 29820 35870 29822 35922
rect 29874 35870 29876 35922
rect 29820 35858 29876 35870
rect 28812 35588 28868 35598
rect 28812 35494 28868 35532
rect 30268 35588 30324 35598
rect 30268 35494 30324 35532
rect 29708 35028 29764 35038
rect 28700 35026 29764 35028
rect 28700 34974 29710 35026
rect 29762 34974 29764 35026
rect 28700 34972 29764 34974
rect 28476 32676 28532 32686
rect 28476 31890 28532 32620
rect 28476 31838 28478 31890
rect 28530 31838 28532 31890
rect 28476 30994 28532 31838
rect 28588 31668 28644 31678
rect 28588 31574 28644 31612
rect 28476 30942 28478 30994
rect 28530 30942 28532 30994
rect 28476 30930 28532 30942
rect 28588 29540 28644 29550
rect 28588 28754 28644 29484
rect 28588 28702 28590 28754
rect 28642 28702 28644 28754
rect 28588 27860 28644 28702
rect 28588 27186 28644 27804
rect 28700 27412 28756 34972
rect 29708 34962 29764 34972
rect 30268 35028 30324 35038
rect 30380 35028 30436 36204
rect 30492 35588 30548 36652
rect 30716 36484 30772 36494
rect 30716 35922 30772 36428
rect 30940 36372 30996 36990
rect 30940 36306 30996 36316
rect 30716 35870 30718 35922
rect 30770 35870 30772 35922
rect 30716 35858 30772 35870
rect 30828 36260 30884 36270
rect 30828 35922 30884 36204
rect 30828 35870 30830 35922
rect 30882 35870 30884 35922
rect 30492 35522 30548 35532
rect 30604 35698 30660 35710
rect 30604 35646 30606 35698
rect 30658 35646 30660 35698
rect 30268 35026 30436 35028
rect 30268 34974 30270 35026
rect 30322 34974 30436 35026
rect 30268 34972 30436 34974
rect 30268 34962 30324 34972
rect 29820 34916 29876 34926
rect 29372 34692 29428 34702
rect 29372 34598 29428 34636
rect 29372 34356 29428 34366
rect 29372 34262 29428 34300
rect 29820 34132 29876 34860
rect 30604 34356 30660 35646
rect 30828 35700 30884 35870
rect 30828 35634 30884 35644
rect 31164 35698 31220 37214
rect 31276 36932 31332 37774
rect 31612 37826 31668 37838
rect 31612 37774 31614 37826
rect 31666 37774 31668 37826
rect 31612 37492 31668 37774
rect 31612 37426 31668 37436
rect 31836 37492 31892 38612
rect 32732 38162 32788 39452
rect 32732 38110 32734 38162
rect 32786 38110 32788 38162
rect 32732 38098 32788 38110
rect 34300 38164 34356 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34412 38164 34468 38174
rect 34300 38162 34468 38164
rect 34300 38110 34414 38162
rect 34466 38110 34468 38162
rect 34300 38108 34468 38110
rect 34412 38098 34468 38108
rect 33740 38050 33796 38062
rect 33740 37998 33742 38050
rect 33794 37998 33796 38050
rect 31836 37426 31892 37436
rect 32396 37492 32452 37502
rect 32396 37398 32452 37436
rect 31388 37380 31444 37390
rect 31388 37286 31444 37324
rect 32732 37380 32788 37390
rect 31500 37268 31556 37278
rect 31500 37174 31556 37212
rect 31276 36866 31332 36876
rect 31948 37154 32004 37166
rect 31948 37102 31950 37154
rect 32002 37102 32004 37154
rect 31948 36708 32004 37102
rect 32732 37156 32788 37324
rect 33740 37380 33796 37998
rect 35420 38052 35476 38062
rect 35420 38050 35588 38052
rect 35420 37998 35422 38050
rect 35474 37998 35588 38050
rect 35420 37996 35588 37998
rect 35420 37986 35476 37996
rect 34972 37492 35028 37502
rect 34972 37398 35028 37436
rect 33740 37314 33796 37324
rect 33628 37268 33684 37278
rect 33292 37156 33348 37166
rect 32732 37100 33124 37156
rect 32508 36932 32564 36942
rect 32396 36876 32508 36932
rect 31948 36652 32228 36708
rect 32060 36484 32116 36494
rect 31948 36372 32004 36382
rect 31948 36278 32004 36316
rect 31948 35924 32004 35934
rect 32060 35924 32116 36428
rect 31948 35922 32116 35924
rect 31948 35870 31950 35922
rect 32002 35870 32116 35922
rect 31948 35868 32116 35870
rect 31948 35858 32004 35868
rect 31164 35646 31166 35698
rect 31218 35646 31220 35698
rect 31164 35634 31220 35646
rect 31836 35698 31892 35710
rect 31836 35646 31838 35698
rect 31890 35646 31892 35698
rect 31836 35026 31892 35646
rect 32060 35700 32116 35710
rect 32060 35606 32116 35644
rect 32172 35476 32228 36652
rect 31836 34974 31838 35026
rect 31890 34974 31892 35026
rect 31836 34962 31892 34974
rect 31948 35420 32228 35476
rect 30828 34916 30884 34926
rect 30716 34356 30772 34366
rect 30604 34354 30772 34356
rect 30604 34302 30718 34354
rect 30770 34302 30772 34354
rect 30604 34300 30772 34302
rect 30716 34290 30772 34300
rect 30828 34356 30884 34860
rect 31388 34916 31444 34926
rect 31388 34822 31444 34860
rect 30940 34692 30996 34702
rect 30940 34598 30996 34636
rect 31612 34692 31668 34702
rect 31836 34692 31892 34702
rect 31612 34690 31780 34692
rect 31612 34638 31614 34690
rect 31666 34638 31780 34690
rect 31612 34636 31780 34638
rect 31612 34626 31668 34636
rect 30828 34262 30884 34300
rect 30940 34300 31444 34356
rect 29820 34020 29876 34076
rect 30492 34132 30548 34142
rect 30492 34038 30548 34076
rect 30604 34130 30660 34142
rect 30604 34078 30606 34130
rect 30658 34078 30660 34130
rect 29708 34018 29876 34020
rect 29708 33966 29822 34018
rect 29874 33966 29876 34018
rect 29708 33964 29876 33966
rect 29148 31780 29204 31790
rect 29148 31686 29204 31724
rect 29260 31668 29316 31678
rect 29260 31574 29316 31612
rect 29260 30884 29316 30894
rect 29148 30212 29204 30222
rect 29148 30118 29204 30156
rect 29260 30210 29316 30828
rect 29260 30158 29262 30210
rect 29314 30158 29316 30210
rect 29260 30146 29316 30158
rect 29596 29876 29652 29886
rect 29708 29876 29764 33964
rect 29820 33954 29876 33964
rect 30604 33908 30660 34078
rect 30940 33908 30996 34300
rect 31388 34242 31444 34300
rect 31388 34190 31390 34242
rect 31442 34190 31444 34242
rect 31388 34178 31444 34190
rect 30604 33852 30996 33908
rect 31052 34130 31108 34142
rect 31052 34078 31054 34130
rect 31106 34078 31108 34130
rect 30380 33684 30436 33694
rect 30380 33346 30436 33628
rect 30380 33294 30382 33346
rect 30434 33294 30436 33346
rect 30380 33282 30436 33294
rect 30492 33236 30548 33246
rect 30492 33142 30548 33180
rect 30716 33124 30772 33134
rect 30716 33122 30996 33124
rect 30716 33070 30718 33122
rect 30770 33070 30996 33122
rect 30716 33068 30996 33070
rect 30716 33058 30772 33068
rect 30828 32788 30884 32798
rect 30828 32694 30884 32732
rect 30604 32676 30660 32686
rect 30604 32674 30772 32676
rect 30604 32622 30606 32674
rect 30658 32622 30772 32674
rect 30604 32620 30772 32622
rect 30604 32610 30660 32620
rect 30492 32562 30548 32574
rect 30492 32510 30494 32562
rect 30546 32510 30548 32562
rect 30492 31892 30548 32510
rect 30492 31826 30548 31836
rect 29820 31668 29876 31678
rect 29820 31574 29876 31612
rect 30604 31668 30660 31678
rect 30604 30772 30660 31612
rect 30716 31444 30772 32620
rect 30940 32340 30996 33068
rect 31052 32674 31108 34078
rect 31724 34020 31780 34636
rect 31836 34598 31892 34636
rect 31724 33964 31892 34020
rect 31612 33458 31668 33470
rect 31612 33406 31614 33458
rect 31666 33406 31668 33458
rect 31052 32622 31054 32674
rect 31106 32622 31108 32674
rect 31052 32610 31108 32622
rect 31500 33348 31556 33358
rect 31388 32450 31444 32462
rect 31388 32398 31390 32450
rect 31442 32398 31444 32450
rect 30940 32284 31332 32340
rect 30940 32116 30996 32126
rect 30828 32060 30940 32116
rect 30828 31666 30884 32060
rect 30940 32050 30996 32060
rect 30940 31892 30996 31902
rect 30940 31798 30996 31836
rect 31276 31778 31332 32284
rect 31388 31892 31444 32398
rect 31500 32116 31556 33292
rect 31500 32050 31556 32060
rect 31388 31826 31444 31836
rect 31276 31726 31278 31778
rect 31330 31726 31332 31778
rect 31276 31714 31332 31726
rect 31500 31668 31556 31678
rect 30828 31614 30830 31666
rect 30882 31614 30884 31666
rect 30828 31602 30884 31614
rect 31388 31666 31556 31668
rect 31388 31614 31502 31666
rect 31554 31614 31556 31666
rect 31388 31612 31556 31614
rect 30716 31378 30772 31388
rect 31164 31444 31220 31454
rect 31388 31444 31444 31612
rect 31500 31602 31556 31612
rect 31612 31668 31668 33406
rect 31836 33460 31892 33964
rect 31948 33684 32004 35420
rect 32396 35252 32452 36876
rect 32508 36866 32564 36876
rect 32732 36706 32788 37100
rect 32732 36654 32734 36706
rect 32786 36654 32788 36706
rect 32732 36642 32788 36654
rect 32844 36932 32900 36942
rect 32844 36482 32900 36876
rect 32844 36430 32846 36482
rect 32898 36430 32900 36482
rect 32844 36418 32900 36430
rect 32508 35698 32564 35710
rect 32508 35646 32510 35698
rect 32562 35646 32564 35698
rect 32508 35588 32564 35646
rect 32956 35698 33012 35710
rect 32956 35646 32958 35698
rect 33010 35646 33012 35698
rect 32956 35588 33012 35646
rect 32508 35532 33012 35588
rect 32396 35196 32676 35252
rect 32508 35028 32564 35038
rect 32172 35026 32564 35028
rect 32172 34974 32510 35026
rect 32562 34974 32564 35026
rect 32172 34972 32564 34974
rect 32060 34914 32116 34926
rect 32060 34862 32062 34914
rect 32114 34862 32116 34914
rect 32060 33908 32116 34862
rect 32172 34018 32228 34972
rect 32508 34962 32564 34972
rect 32396 34802 32452 34814
rect 32396 34750 32398 34802
rect 32450 34750 32452 34802
rect 32172 33966 32174 34018
rect 32226 33966 32228 34018
rect 32172 33954 32228 33966
rect 32284 34130 32340 34142
rect 32284 34078 32286 34130
rect 32338 34078 32340 34130
rect 32060 33842 32116 33852
rect 31948 33628 32228 33684
rect 31948 33460 32004 33470
rect 31836 33458 32004 33460
rect 31836 33406 31950 33458
rect 32002 33406 32004 33458
rect 31836 33404 32004 33406
rect 31948 33394 32004 33404
rect 32172 33348 32228 33628
rect 32172 33282 32228 33292
rect 32284 33236 32340 34078
rect 32396 33684 32452 34750
rect 32396 33618 32452 33628
rect 32508 33908 32564 33918
rect 32508 33460 32564 33852
rect 32508 33394 32564 33404
rect 32284 33142 32340 33180
rect 31724 32562 31780 32574
rect 31724 32510 31726 32562
rect 31778 32510 31780 32562
rect 31724 32004 31780 32510
rect 31724 31938 31780 31948
rect 32508 32004 32564 32014
rect 32060 31892 32116 31902
rect 31836 31780 31892 31790
rect 31836 31686 31892 31724
rect 32060 31778 32116 31836
rect 32060 31726 32062 31778
rect 32114 31726 32116 31778
rect 32060 31714 32116 31726
rect 32508 31778 32564 31948
rect 32508 31726 32510 31778
rect 32562 31726 32564 31778
rect 32508 31714 32564 31726
rect 31612 31602 31668 31612
rect 31724 31554 31780 31566
rect 31724 31502 31726 31554
rect 31778 31502 31780 31554
rect 31220 31388 31444 31444
rect 31500 31444 31556 31454
rect 31164 31378 31220 31388
rect 31500 31106 31556 31388
rect 31612 31220 31668 31230
rect 31612 31126 31668 31164
rect 31500 31054 31502 31106
rect 31554 31054 31556 31106
rect 31500 31042 31556 31054
rect 31724 31108 31780 31502
rect 32284 31554 32340 31566
rect 32284 31502 32286 31554
rect 32338 31502 32340 31554
rect 32172 31108 32228 31118
rect 31724 31052 32172 31108
rect 32172 30994 32228 31052
rect 32172 30942 32174 30994
rect 32226 30942 32228 30994
rect 32172 30930 32228 30942
rect 30604 30706 30660 30716
rect 30716 30882 30772 30894
rect 31276 30884 31332 30894
rect 30716 30830 30718 30882
rect 30770 30830 30772 30882
rect 30604 30098 30660 30110
rect 30604 30046 30606 30098
rect 30658 30046 30660 30098
rect 29652 29820 29764 29876
rect 29820 29986 29876 29998
rect 29820 29934 29822 29986
rect 29874 29934 29876 29986
rect 29596 28754 29652 29820
rect 29596 28702 29598 28754
rect 29650 28702 29652 28754
rect 29596 28690 29652 28702
rect 28700 27346 28756 27356
rect 29148 28644 29204 28654
rect 28588 27134 28590 27186
rect 28642 27134 28644 27186
rect 28588 27122 28644 27134
rect 28364 26226 28420 26236
rect 29036 26852 29092 26862
rect 29036 26290 29092 26796
rect 29036 26238 29038 26290
rect 29090 26238 29092 26290
rect 29036 26226 29092 26238
rect 27580 24670 27582 24722
rect 27634 24670 27636 24722
rect 27580 24658 27636 24670
rect 27692 26180 27748 26190
rect 27132 23998 27134 24050
rect 27186 23998 27188 24050
rect 27132 23986 27188 23998
rect 26684 23828 26740 23838
rect 26796 23828 26852 23838
rect 26740 23826 26964 23828
rect 26740 23774 26798 23826
rect 26850 23774 26964 23826
rect 26740 23772 26964 23774
rect 26684 23762 26740 23772
rect 26796 23734 26852 23772
rect 26684 23268 26740 23278
rect 26572 23266 26740 23268
rect 26572 23214 26686 23266
rect 26738 23214 26740 23266
rect 26572 23212 26740 23214
rect 26460 23156 26516 23166
rect 26460 23062 26516 23100
rect 26572 21700 26628 23212
rect 26684 23202 26740 23212
rect 26796 23154 26852 23166
rect 26796 23102 26798 23154
rect 26850 23102 26852 23154
rect 26796 23044 26852 23102
rect 26796 22978 26852 22988
rect 26908 22484 26964 23772
rect 27020 23716 27076 23726
rect 27020 23714 27188 23716
rect 27020 23662 27022 23714
rect 27074 23662 27188 23714
rect 27020 23660 27188 23662
rect 27020 23650 27076 23660
rect 27132 22708 27188 23660
rect 27244 23714 27300 23726
rect 27244 23662 27246 23714
rect 27298 23662 27300 23714
rect 27244 22932 27300 23662
rect 27356 23714 27412 23726
rect 27356 23662 27358 23714
rect 27410 23662 27412 23714
rect 27356 23378 27412 23662
rect 27356 23326 27358 23378
rect 27410 23326 27412 23378
rect 27356 23314 27412 23326
rect 27692 23268 27748 26124
rect 28476 26178 28532 26190
rect 28476 26126 28478 26178
rect 28530 26126 28532 26178
rect 28252 25284 28308 25294
rect 28140 25282 28308 25284
rect 28140 25230 28254 25282
rect 28306 25230 28308 25282
rect 28140 25228 28308 25230
rect 28140 24948 28196 25228
rect 28252 25218 28308 25228
rect 28140 23716 28196 24892
rect 28252 25060 28308 25070
rect 28252 24722 28308 25004
rect 28476 24836 28532 26126
rect 28812 26178 28868 26190
rect 28812 26126 28814 26178
rect 28866 26126 28868 26178
rect 28812 25508 28868 26126
rect 29148 26180 29204 28588
rect 29820 28644 29876 29934
rect 30380 29986 30436 29998
rect 30380 29934 30382 29986
rect 30434 29934 30436 29986
rect 30380 29316 30436 29934
rect 30380 29250 30436 29260
rect 29820 28578 29876 28588
rect 30380 28644 30436 28654
rect 30380 28550 30436 28588
rect 29708 28084 29764 28094
rect 29708 27990 29764 28028
rect 29596 27860 29652 27870
rect 29596 27298 29652 27804
rect 30380 27860 30436 27870
rect 30380 27766 30436 27804
rect 30604 27748 30660 30046
rect 30716 28756 30772 30830
rect 31164 30882 31332 30884
rect 31164 30830 31278 30882
rect 31330 30830 31332 30882
rect 31164 30828 31332 30830
rect 30940 30210 30996 30222
rect 30940 30158 30942 30210
rect 30994 30158 30996 30210
rect 30716 28690 30772 28700
rect 30828 29652 30884 29662
rect 30716 28084 30772 28094
rect 30716 27990 30772 28028
rect 30828 27970 30884 29596
rect 30940 28084 30996 30158
rect 31052 29986 31108 29998
rect 31052 29934 31054 29986
rect 31106 29934 31108 29986
rect 31052 28866 31108 29934
rect 31052 28814 31054 28866
rect 31106 28814 31108 28866
rect 31052 28802 31108 28814
rect 30940 28018 30996 28028
rect 31052 28532 31108 28542
rect 30828 27918 30830 27970
rect 30882 27918 30884 27970
rect 30828 27906 30884 27918
rect 30604 27682 30660 27692
rect 30716 27300 30772 27310
rect 29596 27246 29598 27298
rect 29650 27246 29652 27298
rect 29596 27234 29652 27246
rect 30380 27298 30772 27300
rect 30380 27246 30718 27298
rect 30770 27246 30772 27298
rect 30380 27244 30772 27246
rect 29820 27188 29876 27198
rect 29484 27076 29540 27086
rect 29260 26964 29316 27002
rect 29260 26898 29316 26908
rect 29484 26908 29540 27020
rect 29820 26962 29876 27132
rect 29820 26910 29822 26962
rect 29874 26910 29876 26962
rect 29484 26852 29652 26908
rect 29820 26898 29876 26910
rect 30380 26962 30436 27244
rect 30716 27234 30772 27244
rect 30380 26910 30382 26962
rect 30434 26910 30436 26962
rect 30380 26898 30436 26910
rect 30940 27074 30996 27086
rect 30940 27022 30942 27074
rect 30994 27022 30996 27074
rect 29484 26290 29540 26302
rect 29484 26238 29486 26290
rect 29538 26238 29540 26290
rect 29148 26114 29204 26124
rect 29260 26178 29316 26190
rect 29260 26126 29262 26178
rect 29314 26126 29316 26178
rect 28812 25442 28868 25452
rect 28476 24770 28532 24780
rect 28588 25282 28644 25294
rect 28588 25230 28590 25282
rect 28642 25230 28644 25282
rect 28252 24670 28254 24722
rect 28306 24670 28308 24722
rect 28252 24658 28308 24670
rect 28588 24724 28644 25230
rect 29260 25060 29316 26126
rect 29484 26180 29540 26238
rect 29484 26114 29540 26124
rect 29596 26068 29652 26852
rect 30940 26852 30996 27022
rect 30940 26786 30996 26796
rect 29596 25506 29652 26012
rect 29596 25454 29598 25506
rect 29650 25454 29652 25506
rect 29596 25442 29652 25454
rect 29708 26290 29764 26302
rect 29708 26238 29710 26290
rect 29762 26238 29764 26290
rect 29708 25284 29764 26238
rect 29932 26292 29988 26302
rect 29988 26236 30100 26292
rect 29932 26226 29988 26236
rect 29820 25508 29876 25518
rect 29820 25506 29988 25508
rect 29820 25454 29822 25506
rect 29874 25454 29988 25506
rect 29820 25452 29988 25454
rect 29820 25442 29876 25452
rect 29820 25284 29876 25294
rect 29708 25282 29876 25284
rect 29708 25230 29822 25282
rect 29874 25230 29876 25282
rect 29708 25228 29876 25230
rect 29820 25218 29876 25228
rect 29260 24994 29316 25004
rect 29372 24836 29428 24846
rect 29596 24836 29652 24846
rect 29428 24780 29540 24836
rect 29372 24770 29428 24780
rect 28476 24162 28532 24174
rect 28476 24110 28478 24162
rect 28530 24110 28532 24162
rect 28252 23938 28308 23950
rect 28252 23886 28254 23938
rect 28306 23886 28308 23938
rect 28252 23828 28308 23886
rect 28364 23940 28420 23950
rect 28364 23846 28420 23884
rect 28252 23762 28308 23772
rect 28140 23650 28196 23660
rect 27748 23212 27972 23268
rect 27692 23202 27748 23212
rect 27916 23154 27972 23212
rect 27916 23102 27918 23154
rect 27970 23102 27972 23154
rect 27692 23044 27748 23054
rect 27692 22950 27748 22988
rect 27244 22866 27300 22876
rect 27132 22652 27860 22708
rect 27132 22484 27188 22494
rect 26908 22482 27188 22484
rect 26908 22430 27134 22482
rect 27186 22430 27188 22482
rect 26908 22428 27188 22430
rect 27132 22418 27188 22428
rect 27468 22148 27524 22158
rect 27468 22054 27524 22092
rect 26572 21634 26628 21644
rect 27580 21700 27636 21710
rect 27804 21700 27860 22652
rect 27916 22482 27972 23102
rect 27916 22430 27918 22482
rect 27970 22430 27972 22482
rect 27916 22418 27972 22430
rect 28476 22484 28532 24110
rect 28588 23548 28644 24668
rect 29484 24050 29540 24780
rect 29596 24162 29652 24780
rect 29596 24110 29598 24162
rect 29650 24110 29652 24162
rect 29596 24098 29652 24110
rect 29484 23998 29486 24050
rect 29538 23998 29540 24050
rect 29484 23604 29540 23998
rect 28588 23492 28980 23548
rect 29484 23538 29540 23548
rect 28588 23154 28644 23166
rect 28588 23102 28590 23154
rect 28642 23102 28644 23154
rect 28588 22596 28644 23102
rect 28700 23044 28756 23054
rect 28700 22950 28756 22988
rect 28588 22502 28644 22540
rect 28476 22418 28532 22428
rect 28476 22258 28532 22270
rect 28476 22206 28478 22258
rect 28530 22206 28532 22258
rect 27916 21700 27972 21710
rect 27804 21698 27972 21700
rect 27804 21646 27918 21698
rect 27970 21646 27972 21698
rect 27804 21644 27972 21646
rect 26908 21588 26964 21598
rect 26908 21494 26964 21532
rect 26684 21028 26740 21038
rect 26684 20914 26740 20972
rect 27580 21026 27636 21644
rect 27916 21634 27972 21644
rect 28476 21700 28532 22206
rect 28476 21634 28532 21644
rect 27580 20974 27582 21026
rect 27634 20974 27636 21026
rect 27580 20962 27636 20974
rect 28364 21588 28420 21598
rect 26684 20862 26686 20914
rect 26738 20862 26740 20914
rect 26684 20850 26740 20862
rect 27692 20804 27748 20814
rect 27692 20710 27748 20748
rect 27356 20690 27412 20702
rect 27356 20638 27358 20690
rect 27410 20638 27412 20690
rect 26572 20132 26628 20142
rect 26572 20020 26628 20076
rect 26460 20018 26628 20020
rect 26460 19966 26574 20018
rect 26626 19966 26628 20018
rect 26460 19964 26628 19966
rect 26460 19684 26516 19964
rect 26572 19954 26628 19964
rect 26684 20020 26740 20030
rect 26684 19926 26740 19964
rect 26796 20018 26852 20030
rect 26796 19966 26798 20018
rect 26850 19966 26852 20018
rect 26460 19618 26516 19628
rect 26572 19796 26628 19806
rect 26348 19182 26350 19234
rect 26402 19182 26404 19234
rect 26236 19124 26292 19134
rect 26236 19030 26292 19068
rect 25788 18386 25844 18396
rect 25564 18284 25732 18340
rect 25676 18228 25732 18284
rect 25900 18338 25956 18350
rect 25900 18286 25902 18338
rect 25954 18286 25956 18338
rect 25900 18228 25956 18286
rect 25676 18172 25956 18228
rect 25900 17780 25956 18172
rect 26348 18340 26404 19182
rect 26572 19122 26628 19740
rect 26572 19070 26574 19122
rect 26626 19070 26628 19122
rect 26572 19058 26628 19070
rect 26348 17892 26404 18284
rect 26348 17826 26404 17836
rect 26796 18452 26852 19966
rect 27244 20018 27300 20030
rect 27244 19966 27246 20018
rect 27298 19966 27300 20018
rect 27244 19908 27300 19966
rect 27244 19842 27300 19852
rect 27356 18788 27412 20638
rect 28140 20578 28196 20590
rect 28140 20526 28142 20578
rect 28194 20526 28196 20578
rect 26796 18338 26852 18396
rect 26908 18732 27412 18788
rect 27580 19906 27636 19918
rect 28028 19908 28084 19918
rect 28140 19908 28196 20526
rect 28364 19908 28420 21532
rect 28812 21474 28868 21486
rect 28812 21422 28814 21474
rect 28866 21422 28868 21474
rect 28812 20692 28868 21422
rect 28924 21252 28980 23492
rect 29932 23492 29988 25452
rect 30044 25506 30100 26236
rect 30380 26180 30436 26190
rect 30380 25620 30436 26124
rect 30044 25454 30046 25506
rect 30098 25454 30100 25506
rect 30044 25442 30100 25454
rect 30156 25564 30436 25620
rect 30716 26178 30772 26190
rect 30716 26126 30718 26178
rect 30770 26126 30772 26178
rect 30716 25620 30772 26126
rect 30156 25172 30212 25564
rect 30716 25554 30772 25564
rect 30828 25508 30884 25518
rect 30268 25396 30324 25406
rect 30268 25302 30324 25340
rect 30156 25116 30436 25172
rect 30380 23940 30436 25116
rect 30492 24836 30548 24846
rect 30492 24742 30548 24780
rect 30380 23846 30436 23884
rect 30492 23828 30548 23838
rect 30828 23828 30884 25452
rect 30548 23772 30884 23828
rect 30268 23716 30324 23726
rect 29932 23436 30100 23492
rect 29708 23380 29764 23390
rect 29036 22932 29092 22942
rect 29036 22370 29092 22876
rect 29484 22596 29540 22606
rect 29484 22502 29540 22540
rect 29708 22594 29764 23324
rect 29708 22542 29710 22594
rect 29762 22542 29764 22594
rect 29708 22530 29764 22542
rect 29932 23044 29988 23054
rect 29932 22594 29988 22988
rect 29932 22542 29934 22594
rect 29986 22542 29988 22594
rect 29932 22530 29988 22542
rect 29036 22318 29038 22370
rect 29090 22318 29092 22370
rect 29036 22306 29092 22318
rect 30044 21812 30100 23436
rect 30156 22484 30212 22494
rect 30156 22390 30212 22428
rect 30268 21812 30324 23660
rect 30044 21746 30100 21756
rect 30156 21756 30324 21812
rect 29260 21700 29316 21710
rect 29260 21606 29316 21644
rect 29708 21588 29764 21598
rect 29764 21532 29876 21588
rect 29708 21494 29764 21532
rect 28924 21186 28980 21196
rect 29260 21028 29316 21038
rect 29260 20934 29316 20972
rect 29820 20914 29876 21532
rect 29820 20862 29822 20914
rect 29874 20862 29876 20914
rect 29820 20850 29876 20862
rect 30156 21586 30212 21756
rect 30156 21534 30158 21586
rect 30210 21534 30212 21586
rect 30156 20804 30212 21534
rect 30156 20738 30212 20748
rect 30268 21588 30324 21598
rect 30492 21588 30548 23772
rect 30604 23604 30660 23614
rect 30604 22482 30660 23548
rect 30604 22430 30606 22482
rect 30658 22430 30660 22482
rect 30604 22418 30660 22430
rect 31052 22372 31108 28476
rect 31164 27860 31220 30828
rect 31276 30818 31332 30828
rect 32060 30884 32116 30894
rect 32060 30790 32116 30828
rect 31948 30772 32004 30782
rect 31276 30212 31332 30222
rect 31276 30118 31332 30156
rect 31948 30098 32004 30716
rect 32284 30436 32340 31502
rect 32396 30996 32452 31006
rect 32396 30902 32452 30940
rect 32284 30370 32340 30380
rect 32508 30770 32564 30782
rect 32508 30718 32510 30770
rect 32562 30718 32564 30770
rect 31948 30046 31950 30098
rect 32002 30046 32004 30098
rect 31948 30034 32004 30046
rect 32396 30212 32452 30222
rect 32060 29652 32116 29662
rect 32060 29558 32116 29596
rect 31388 29540 31444 29550
rect 31388 29446 31444 29484
rect 31724 29316 31780 29326
rect 31500 28756 31556 28766
rect 31500 28662 31556 28700
rect 31276 28644 31332 28654
rect 31276 28642 31444 28644
rect 31276 28590 31278 28642
rect 31330 28590 31444 28642
rect 31276 28588 31444 28590
rect 31276 28578 31332 28588
rect 31388 27972 31444 28588
rect 31724 28642 31780 29260
rect 31724 28590 31726 28642
rect 31778 28590 31780 28642
rect 31724 28532 31780 28590
rect 31948 28644 32004 28654
rect 32172 28644 32228 28654
rect 31948 28642 32172 28644
rect 31948 28590 31950 28642
rect 32002 28590 32172 28642
rect 31948 28588 32172 28590
rect 31948 28578 32004 28588
rect 32172 28578 32228 28588
rect 32396 28532 32452 30156
rect 32508 30100 32564 30718
rect 32508 30034 32564 30044
rect 32508 29652 32564 29662
rect 32620 29652 32676 35196
rect 32732 34804 32788 34814
rect 32732 34802 32900 34804
rect 32732 34750 32734 34802
rect 32786 34750 32900 34802
rect 32732 34748 32900 34750
rect 32732 34738 32788 34748
rect 32732 33572 32788 33582
rect 32732 33346 32788 33516
rect 32732 33294 32734 33346
rect 32786 33294 32788 33346
rect 32732 33282 32788 33294
rect 32732 32788 32788 32798
rect 32844 32788 32900 34748
rect 32788 32732 32900 32788
rect 32956 34802 33012 34814
rect 32956 34750 32958 34802
rect 33010 34750 33012 34802
rect 32956 33348 33012 34750
rect 33068 33572 33124 37100
rect 33292 37154 33572 37156
rect 33292 37102 33294 37154
rect 33346 37102 33572 37154
rect 33292 37100 33572 37102
rect 33292 37090 33348 37100
rect 33516 36932 33572 37100
rect 33628 37044 33684 37212
rect 34076 37156 34132 37166
rect 34524 37156 34580 37166
rect 34076 37154 34580 37156
rect 34076 37102 34078 37154
rect 34130 37102 34526 37154
rect 34578 37102 34580 37154
rect 34076 37100 34580 37102
rect 33628 36988 33908 37044
rect 33516 36876 33684 36932
rect 33180 36708 33236 36718
rect 33180 35924 33236 36652
rect 33404 36484 33460 36494
rect 33404 36390 33460 36428
rect 33180 35922 33460 35924
rect 33180 35870 33182 35922
rect 33234 35870 33460 35922
rect 33180 35868 33460 35870
rect 33180 35858 33236 35868
rect 33292 35698 33348 35710
rect 33292 35646 33294 35698
rect 33346 35646 33348 35698
rect 33292 35476 33348 35646
rect 33292 35410 33348 35420
rect 33404 35026 33460 35868
rect 33628 35588 33684 36876
rect 33740 35700 33796 35710
rect 33740 35606 33796 35644
rect 33628 35522 33684 35532
rect 33852 35476 33908 36988
rect 34076 36932 34132 37100
rect 34524 37090 34580 37100
rect 34076 36866 34132 36876
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35532 36708 35588 37996
rect 35532 36642 35588 36652
rect 36540 36708 36596 36718
rect 36540 36614 36596 36652
rect 34412 36260 34468 36270
rect 34412 35922 34468 36204
rect 35756 36260 35812 36270
rect 35756 36166 35812 36204
rect 34412 35870 34414 35922
rect 34466 35870 34468 35922
rect 34412 35858 34468 35870
rect 33852 35410 33908 35420
rect 34300 35588 34356 35598
rect 33404 34974 33406 35026
rect 33458 34974 33460 35026
rect 33404 34962 33460 34974
rect 33964 34916 34020 34926
rect 33964 34822 34020 34860
rect 33516 34690 33572 34702
rect 33516 34638 33518 34690
rect 33570 34638 33572 34690
rect 33516 34132 33572 34638
rect 34300 34692 34356 35532
rect 34860 35586 34916 35598
rect 34860 35534 34862 35586
rect 34914 35534 34916 35586
rect 34860 35476 34916 35534
rect 34860 35410 34916 35420
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34412 34692 34468 34702
rect 34300 34690 34468 34692
rect 34300 34638 34414 34690
rect 34466 34638 34468 34690
rect 34300 34636 34468 34638
rect 33628 34132 33684 34142
rect 33516 34076 33628 34132
rect 33628 34038 33684 34076
rect 33292 34018 33348 34030
rect 33292 33966 33294 34018
rect 33346 33966 33348 34018
rect 33292 33684 33348 33966
rect 34076 34018 34132 34030
rect 34076 33966 34078 34018
rect 34130 33966 34132 34018
rect 33740 33684 33796 33694
rect 34076 33684 34132 33966
rect 33292 33628 33572 33684
rect 33124 33516 33460 33572
rect 33068 33506 33124 33516
rect 32732 32722 32788 32732
rect 32956 32562 33012 33292
rect 32956 32510 32958 32562
rect 33010 32510 33012 32562
rect 32956 32498 33012 32510
rect 33180 33346 33236 33358
rect 33180 33294 33182 33346
rect 33234 33294 33236 33346
rect 33180 32564 33236 33294
rect 33404 32786 33460 33516
rect 33516 33236 33572 33628
rect 33796 33628 34132 33684
rect 33628 33460 33684 33498
rect 33628 33394 33684 33404
rect 33740 33346 33796 33628
rect 33740 33294 33742 33346
rect 33794 33294 33796 33346
rect 33740 33282 33796 33294
rect 34188 33346 34244 33358
rect 34188 33294 34190 33346
rect 34242 33294 34244 33346
rect 33628 33236 33684 33246
rect 33516 33180 33628 33236
rect 33628 33170 33684 33180
rect 33404 32734 33406 32786
rect 33458 32734 33460 32786
rect 33404 32676 33460 32734
rect 34188 32788 34244 33294
rect 34188 32722 34244 32732
rect 33404 32610 33460 32620
rect 34076 32676 34132 32686
rect 34076 32582 34132 32620
rect 33180 32004 33236 32508
rect 33628 32564 33684 32574
rect 33628 32470 33684 32508
rect 33852 32562 33908 32574
rect 33852 32510 33854 32562
rect 33906 32510 33908 32562
rect 33180 31890 33236 31948
rect 33180 31838 33182 31890
rect 33234 31838 33236 31890
rect 33180 31826 33236 31838
rect 33516 32450 33572 32462
rect 33516 32398 33518 32450
rect 33570 32398 33572 32450
rect 33516 31780 33572 32398
rect 33740 31780 33796 31790
rect 33516 31778 33796 31780
rect 33516 31726 33742 31778
rect 33794 31726 33796 31778
rect 33516 31724 33796 31726
rect 33740 31714 33796 31724
rect 32732 31668 32788 31678
rect 32732 31666 32900 31668
rect 32732 31614 32734 31666
rect 32786 31614 32900 31666
rect 32732 31612 32900 31614
rect 32732 31602 32788 31612
rect 32508 29650 32676 29652
rect 32508 29598 32510 29650
rect 32562 29598 32676 29650
rect 32508 29596 32676 29598
rect 32508 29540 32564 29596
rect 32508 29474 32564 29484
rect 32508 29092 32564 29102
rect 32508 28866 32564 29036
rect 32508 28814 32510 28866
rect 32562 28814 32564 28866
rect 32508 28802 32564 28814
rect 31724 28466 31780 28476
rect 32284 28530 32452 28532
rect 32284 28478 32398 28530
rect 32450 28478 32452 28530
rect 32284 28476 32452 28478
rect 31836 28418 31892 28430
rect 31836 28366 31838 28418
rect 31890 28366 31892 28418
rect 31388 27916 31780 27972
rect 31164 27794 31220 27804
rect 31500 27748 31556 27758
rect 31500 27654 31556 27692
rect 31500 27298 31556 27310
rect 31500 27246 31502 27298
rect 31554 27246 31556 27298
rect 31500 27076 31556 27246
rect 31724 27298 31780 27916
rect 31724 27246 31726 27298
rect 31778 27246 31780 27298
rect 31724 27234 31780 27246
rect 31836 27076 31892 28366
rect 32284 27972 32340 28476
rect 32396 28466 32452 28476
rect 32508 28532 32564 28542
rect 32508 28438 32564 28476
rect 32396 28084 32452 28094
rect 32452 28028 32564 28084
rect 32396 28018 32452 28028
rect 32060 27916 32340 27972
rect 31500 27020 31892 27076
rect 31948 27860 32004 27870
rect 31948 27188 32004 27804
rect 31948 26908 32004 27132
rect 31388 26852 31444 26862
rect 31276 26850 31444 26852
rect 31276 26798 31390 26850
rect 31442 26798 31444 26850
rect 31276 26796 31444 26798
rect 31164 26292 31220 26302
rect 31164 26198 31220 26236
rect 31276 25508 31332 26796
rect 31388 26786 31444 26796
rect 31836 26852 32004 26908
rect 32060 26908 32116 27916
rect 32172 27748 32228 27758
rect 32172 27074 32228 27692
rect 32284 27746 32340 27758
rect 32284 27694 32286 27746
rect 32338 27694 32340 27746
rect 32284 27636 32340 27694
rect 32284 27570 32340 27580
rect 32172 27022 32174 27074
rect 32226 27022 32228 27074
rect 32172 27010 32228 27022
rect 32508 27074 32564 28028
rect 32620 27860 32676 29596
rect 32844 31220 32900 31612
rect 33404 31666 33460 31678
rect 33404 31614 33406 31666
rect 33458 31614 33460 31666
rect 32620 27794 32676 27804
rect 32732 29204 32788 29214
rect 32732 27636 32788 29148
rect 32844 28980 32900 31164
rect 33068 31556 33124 31566
rect 33068 31218 33124 31500
rect 33068 31166 33070 31218
rect 33122 31166 33124 31218
rect 33068 30884 33124 31166
rect 33292 31108 33348 31118
rect 33292 31014 33348 31052
rect 33068 30818 33124 30828
rect 33180 30882 33236 30894
rect 33180 30830 33182 30882
rect 33234 30830 33236 30882
rect 33180 30212 33236 30830
rect 33404 30324 33460 31614
rect 33852 31666 33908 32510
rect 34188 32564 34244 32574
rect 34188 32470 34244 32508
rect 33852 31614 33854 31666
rect 33906 31614 33908 31666
rect 33852 31602 33908 31614
rect 34076 31556 34132 31566
rect 34076 31462 34132 31500
rect 33404 30258 33460 30268
rect 33516 31444 33572 31454
rect 33180 30146 33236 30156
rect 33516 30210 33572 31388
rect 33740 30996 33796 31006
rect 33740 30902 33796 30940
rect 33516 30158 33518 30210
rect 33570 30158 33572 30210
rect 33516 30146 33572 30158
rect 33964 29986 34020 29998
rect 33964 29934 33966 29986
rect 34018 29934 34020 29986
rect 33516 29426 33572 29438
rect 33516 29374 33518 29426
rect 33570 29374 33572 29426
rect 33068 29314 33124 29326
rect 33068 29262 33070 29314
rect 33122 29262 33124 29314
rect 32956 28980 33012 28990
rect 32844 28924 32956 28980
rect 32956 28914 33012 28924
rect 33068 28644 33124 29262
rect 33516 29204 33572 29374
rect 33964 29428 34020 29934
rect 34412 29652 34468 34636
rect 35084 34132 35140 34142
rect 35084 33572 35140 34076
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35084 33516 35364 33572
rect 35084 33348 35140 33358
rect 35084 33254 35140 33292
rect 35308 33346 35364 33516
rect 35308 33294 35310 33346
rect 35362 33294 35364 33346
rect 35308 33282 35364 33294
rect 34972 33236 35028 33246
rect 34860 30996 34916 31006
rect 34412 29586 34468 29596
rect 34524 30100 34580 30110
rect 34524 29650 34580 30044
rect 34524 29598 34526 29650
rect 34578 29598 34580 29650
rect 34524 29586 34580 29598
rect 33964 29334 34020 29372
rect 34748 29426 34804 29438
rect 34748 29374 34750 29426
rect 34802 29374 34804 29426
rect 33516 29138 33572 29148
rect 34636 29314 34692 29326
rect 34636 29262 34638 29314
rect 34690 29262 34692 29314
rect 33292 28980 33348 28990
rect 33068 28578 33124 28588
rect 33180 28756 33236 28766
rect 32956 28084 33012 28094
rect 32956 27990 33012 28028
rect 33180 28082 33236 28700
rect 33180 28030 33182 28082
rect 33234 28030 33236 28082
rect 33180 28018 33236 28030
rect 33292 27970 33348 28924
rect 33964 28756 34020 28766
rect 33964 28662 34020 28700
rect 33516 28642 33572 28654
rect 33516 28590 33518 28642
rect 33570 28590 33572 28642
rect 33404 28532 33460 28542
rect 33404 28438 33460 28476
rect 33292 27918 33294 27970
rect 33346 27918 33348 27970
rect 33292 27906 33348 27918
rect 32732 27570 32788 27580
rect 33180 27860 33236 27870
rect 32508 27022 32510 27074
rect 32562 27022 32564 27074
rect 32508 27010 32564 27022
rect 32284 26962 32340 26974
rect 32284 26910 32286 26962
rect 32338 26910 32340 26962
rect 32284 26908 32340 26910
rect 32060 26852 32340 26908
rect 31612 26178 31668 26190
rect 31612 26126 31614 26178
rect 31666 26126 31668 26178
rect 31612 26068 31668 26126
rect 31612 26002 31668 26012
rect 31276 25442 31332 25452
rect 31500 25508 31556 25518
rect 31556 25452 31668 25508
rect 31500 25414 31556 25452
rect 31164 25396 31220 25406
rect 31164 24948 31220 25340
rect 31164 24892 31556 24948
rect 31500 24834 31556 24892
rect 31500 24782 31502 24834
rect 31554 24782 31556 24834
rect 31500 24770 31556 24782
rect 31276 24612 31332 24622
rect 31612 24612 31668 25452
rect 31724 25394 31780 25406
rect 31724 25342 31726 25394
rect 31778 25342 31780 25394
rect 31724 24836 31780 25342
rect 31724 24722 31780 24780
rect 31724 24670 31726 24722
rect 31778 24670 31780 24722
rect 31724 24658 31780 24670
rect 31276 24610 31668 24612
rect 31276 24558 31278 24610
rect 31330 24558 31668 24610
rect 31276 24556 31668 24558
rect 31276 24546 31332 24556
rect 31836 24164 31892 26852
rect 33068 26850 33124 26862
rect 33068 26798 33070 26850
rect 33122 26798 33124 26850
rect 31948 26740 32004 26750
rect 33068 26740 33124 26798
rect 31948 26402 32004 26684
rect 31948 26350 31950 26402
rect 32002 26350 32004 26402
rect 31948 26338 32004 26350
rect 32396 26684 33124 26740
rect 32172 26290 32228 26302
rect 32172 26238 32174 26290
rect 32226 26238 32228 26290
rect 32060 26178 32116 26190
rect 32060 26126 32062 26178
rect 32114 26126 32116 26178
rect 32060 25844 32116 26126
rect 32060 25778 32116 25788
rect 31724 24108 31892 24164
rect 31948 25732 32004 25742
rect 31164 23714 31220 23726
rect 31164 23662 31166 23714
rect 31218 23662 31220 23714
rect 31164 23044 31220 23662
rect 31724 23380 31780 24108
rect 31724 23324 31892 23380
rect 31164 22950 31220 22988
rect 31388 23154 31444 23166
rect 31388 23102 31390 23154
rect 31442 23102 31444 23154
rect 31388 22484 31444 23102
rect 31388 22418 31444 22428
rect 31612 22484 31668 22494
rect 31612 22390 31668 22428
rect 31052 22316 31332 22372
rect 31052 22146 31108 22158
rect 31052 22094 31054 22146
rect 31106 22094 31108 22146
rect 30940 21812 30996 21822
rect 30940 21718 30996 21756
rect 30324 21532 30548 21588
rect 30604 21586 30660 21598
rect 30604 21534 30606 21586
rect 30658 21534 30660 21586
rect 29148 20692 29204 20702
rect 28812 20690 29204 20692
rect 28812 20638 29150 20690
rect 29202 20638 29204 20690
rect 28812 20636 29204 20638
rect 28588 20580 28644 20590
rect 28588 20486 28644 20524
rect 29148 20132 29204 20636
rect 29260 20580 29316 20590
rect 29260 20486 29316 20524
rect 30268 20578 30324 21532
rect 30604 21028 30660 21534
rect 30828 21588 30884 21598
rect 31052 21588 31108 22094
rect 30884 21532 31108 21588
rect 31164 21586 31220 21598
rect 31164 21534 31166 21586
rect 31218 21534 31220 21586
rect 30828 21494 30884 21532
rect 31164 21028 31220 21534
rect 30604 20962 30660 20972
rect 30940 20972 31220 21028
rect 30940 20916 30996 20972
rect 30268 20526 30270 20578
rect 30322 20526 30324 20578
rect 29148 20038 29204 20076
rect 29260 20020 29316 20030
rect 30268 20020 30324 20526
rect 30716 20914 30996 20916
rect 30716 20862 30942 20914
rect 30994 20862 30996 20914
rect 30716 20860 30996 20862
rect 30604 20244 30660 20254
rect 30716 20244 30772 20860
rect 30940 20850 30996 20860
rect 30604 20242 30772 20244
rect 30604 20190 30606 20242
rect 30658 20190 30772 20242
rect 30604 20188 30772 20190
rect 31164 20802 31220 20814
rect 31164 20750 31166 20802
rect 31218 20750 31220 20802
rect 30604 20178 30660 20188
rect 30380 20020 30436 20030
rect 30268 19964 30380 20020
rect 28476 19908 28532 19918
rect 27580 19854 27582 19906
rect 27634 19854 27636 19906
rect 26908 18450 26964 18732
rect 26908 18398 26910 18450
rect 26962 18398 26964 18450
rect 26908 18386 26964 18398
rect 26796 18286 26798 18338
rect 26850 18286 26852 18338
rect 25900 17714 25956 17724
rect 25228 17444 25284 17454
rect 25228 17108 25284 17388
rect 25228 16882 25284 17052
rect 25228 16830 25230 16882
rect 25282 16830 25284 16882
rect 25228 16818 25284 16830
rect 25452 16098 25508 17612
rect 26684 17444 26740 17454
rect 26124 16996 26180 17006
rect 25452 16046 25454 16098
rect 25506 16046 25508 16098
rect 25452 16034 25508 16046
rect 25900 16772 25956 16782
rect 25116 15988 25172 15998
rect 25116 15986 25396 15988
rect 25116 15934 25118 15986
rect 25170 15934 25396 15986
rect 25116 15932 25396 15934
rect 25116 15922 25172 15932
rect 24668 15474 24724 15484
rect 24108 15426 24164 15438
rect 24108 15374 24110 15426
rect 24162 15374 24164 15426
rect 23212 14354 23268 14364
rect 23324 15092 23492 15148
rect 23772 15314 23828 15326
rect 23772 15262 23774 15314
rect 23826 15262 23828 15314
rect 22876 13022 22878 13074
rect 22930 13022 22932 13074
rect 22876 12964 22932 13022
rect 22876 12898 22932 12908
rect 22988 12292 23044 12302
rect 22988 12198 23044 12236
rect 22764 11974 22820 12012
rect 23100 12178 23156 12190
rect 23100 12126 23102 12178
rect 23154 12126 23156 12178
rect 22652 11454 22654 11506
rect 22706 11454 22708 11506
rect 22652 11442 22708 11454
rect 22876 11956 22932 11966
rect 22428 9774 22430 9826
rect 22482 9774 22484 9826
rect 22428 9716 22484 9774
rect 22876 11394 22932 11900
rect 22876 11342 22878 11394
rect 22930 11342 22932 11394
rect 22876 10500 22932 11342
rect 22484 9660 22708 9716
rect 22428 9650 22484 9660
rect 21868 9266 22484 9268
rect 21868 9214 21870 9266
rect 21922 9214 22484 9266
rect 21868 9212 22484 9214
rect 21868 9202 21924 9212
rect 22428 9042 22484 9212
rect 22652 9044 22708 9660
rect 22428 8990 22430 9042
rect 22482 8990 22484 9042
rect 22428 8978 22484 8990
rect 22540 9042 22708 9044
rect 22540 8990 22654 9042
rect 22706 8990 22708 9042
rect 22540 8988 22708 8990
rect 21420 8318 21422 8370
rect 21474 8318 21476 8370
rect 21308 7698 21364 7710
rect 21308 7646 21310 7698
rect 21362 7646 21364 7698
rect 21308 6914 21364 7646
rect 21308 6862 21310 6914
rect 21362 6862 21364 6914
rect 21308 6850 21364 6862
rect 21420 6804 21476 8318
rect 22204 8258 22260 8270
rect 22204 8206 22206 8258
rect 22258 8206 22260 8258
rect 21420 6802 21812 6804
rect 21420 6750 21422 6802
rect 21474 6750 21812 6802
rect 21420 6748 21812 6750
rect 21420 6738 21476 6748
rect 21756 6692 21812 6748
rect 21980 6692 22036 6702
rect 22204 6692 22260 8206
rect 22316 7700 22372 7710
rect 22540 7700 22596 8988
rect 22652 8978 22708 8988
rect 22876 9042 22932 10444
rect 23100 11844 23156 12126
rect 23100 9725 23156 11788
rect 23100 9673 23102 9725
rect 23154 9673 23156 9725
rect 23100 9661 23156 9673
rect 23212 9716 23268 9726
rect 23212 9266 23268 9660
rect 23212 9214 23214 9266
rect 23266 9214 23268 9266
rect 23212 9202 23268 9214
rect 22876 8990 22878 9042
rect 22930 8990 22932 9042
rect 22876 8978 22932 8990
rect 22316 7698 22596 7700
rect 22316 7646 22318 7698
rect 22370 7646 22596 7698
rect 22316 7644 22596 7646
rect 22652 8258 22708 8270
rect 22652 8206 22654 8258
rect 22706 8206 22708 8258
rect 22316 7634 22372 7644
rect 22652 7588 22708 8206
rect 22652 7522 22708 7532
rect 21756 6690 22148 6692
rect 21756 6638 21982 6690
rect 22034 6638 22148 6690
rect 21756 6636 22148 6638
rect 21980 6626 22036 6636
rect 22092 6468 22148 6636
rect 22204 6626 22260 6636
rect 22428 6468 22484 6478
rect 22092 6412 22428 6468
rect 22428 6374 22484 6412
rect 22204 3668 22260 3678
rect 18396 3378 18452 3388
rect 21084 3378 21140 3388
rect 21532 3666 22260 3668
rect 21532 3614 22206 3666
rect 22258 3614 22260 3666
rect 21532 3612 22260 3614
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 21532 800 21588 3612
rect 22204 3602 22260 3612
rect 23100 3556 23156 3566
rect 21756 3444 21812 3482
rect 23100 3388 23156 3500
rect 21756 3378 21812 3388
rect 22876 3332 23156 3388
rect 23324 3442 23380 15092
rect 23772 13860 23828 15262
rect 23996 14530 24052 14542
rect 23996 14478 23998 14530
rect 24050 14478 24052 14530
rect 23996 14420 24052 14478
rect 24108 14532 24164 15374
rect 25340 15316 25396 15932
rect 25788 15540 25844 15550
rect 25788 15446 25844 15484
rect 25900 15538 25956 16716
rect 25900 15486 25902 15538
rect 25954 15486 25956 15538
rect 25900 15474 25956 15486
rect 26012 16770 26068 16782
rect 26012 16718 26014 16770
rect 26066 16718 26068 16770
rect 26012 15988 26068 16718
rect 25676 15316 25732 15326
rect 26012 15316 26068 15932
rect 25396 15260 25620 15316
rect 25340 15222 25396 15260
rect 24444 15202 24500 15214
rect 24444 15150 24446 15202
rect 24498 15150 24500 15202
rect 24332 14532 24388 14542
rect 24108 14530 24388 14532
rect 24108 14478 24334 14530
rect 24386 14478 24388 14530
rect 24108 14476 24388 14478
rect 23996 14354 24052 14364
rect 24220 14306 24276 14318
rect 24220 14254 24222 14306
rect 24274 14254 24276 14306
rect 24108 13972 24164 13982
rect 24108 13878 24164 13916
rect 23772 13188 23828 13804
rect 23772 13122 23828 13132
rect 23884 13636 23940 13646
rect 23660 12964 23716 12974
rect 23884 12964 23940 13580
rect 24220 13524 24276 14254
rect 24332 13636 24388 14476
rect 24332 13570 24388 13580
rect 24220 13458 24276 13468
rect 23660 12962 23940 12964
rect 23660 12910 23662 12962
rect 23714 12910 23940 12962
rect 23660 12908 23940 12910
rect 23660 11956 23716 12908
rect 23660 11890 23716 11900
rect 23772 12292 23828 12302
rect 23772 11394 23828 12236
rect 23772 11342 23774 11394
rect 23826 11342 23828 11394
rect 23772 10724 23828 11342
rect 24444 11284 24500 15150
rect 25228 15202 25284 15214
rect 25228 15150 25230 15202
rect 25282 15150 25284 15202
rect 24780 14532 24836 14542
rect 24780 14418 24836 14476
rect 24780 14366 24782 14418
rect 24834 14366 24836 14418
rect 24780 13076 24836 14366
rect 25228 14196 25284 15150
rect 25228 14130 25284 14140
rect 25340 15090 25396 15102
rect 25340 15038 25342 15090
rect 25394 15038 25396 15090
rect 25340 13860 25396 15038
rect 25564 13972 25620 15260
rect 25676 15314 26068 15316
rect 25676 15262 25678 15314
rect 25730 15262 26068 15314
rect 25676 15260 26068 15262
rect 26124 16210 26180 16940
rect 26572 16996 26628 17006
rect 26684 16996 26740 17388
rect 26628 16940 26740 16996
rect 26572 16930 26628 16940
rect 26684 16772 26740 16940
rect 26796 16996 26852 18286
rect 26908 17442 26964 17454
rect 26908 17390 26910 17442
rect 26962 17390 26964 17442
rect 26908 17106 26964 17390
rect 26908 17054 26910 17106
rect 26962 17054 26964 17106
rect 26908 17042 26964 17054
rect 26796 16930 26852 16940
rect 26796 16772 26852 16782
rect 26684 16770 26852 16772
rect 26684 16718 26798 16770
rect 26850 16718 26852 16770
rect 26684 16716 26852 16718
rect 26796 16706 26852 16716
rect 27020 16772 27076 18732
rect 27356 18340 27412 18350
rect 27356 18246 27412 18284
rect 27580 18340 27636 19854
rect 27916 19906 28532 19908
rect 27916 19854 28030 19906
rect 28082 19854 28478 19906
rect 28530 19854 28532 19906
rect 27916 19852 28532 19854
rect 27580 18274 27636 18284
rect 27804 18340 27860 18350
rect 27916 18340 27972 19852
rect 28028 19842 28084 19852
rect 28476 19842 28532 19852
rect 28476 19236 28532 19246
rect 28476 19142 28532 19180
rect 27804 18338 27972 18340
rect 27804 18286 27806 18338
rect 27858 18286 27972 18338
rect 27804 18284 27972 18286
rect 28028 19010 28084 19022
rect 28028 18958 28030 19010
rect 28082 18958 28084 19010
rect 27692 17444 27748 17454
rect 27020 16706 27076 16716
rect 27132 17442 27748 17444
rect 27132 17390 27694 17442
rect 27746 17390 27748 17442
rect 27132 17388 27748 17390
rect 26124 16158 26126 16210
rect 26178 16158 26180 16210
rect 25676 15204 25732 15260
rect 25676 15138 25732 15148
rect 26124 14868 26180 16158
rect 26684 16100 26740 16110
rect 26348 15876 26404 15886
rect 26348 15314 26404 15820
rect 26348 15262 26350 15314
rect 26402 15262 26404 15314
rect 26348 15250 26404 15262
rect 26684 15314 26740 16044
rect 27132 15986 27188 17388
rect 27692 17378 27748 17388
rect 27804 16996 27860 18284
rect 28028 18226 28084 18958
rect 29260 19010 29316 19964
rect 30380 19926 30436 19964
rect 29708 19794 29764 19806
rect 29708 19742 29710 19794
rect 29762 19742 29764 19794
rect 29708 19684 29764 19742
rect 29932 19796 29988 19806
rect 29932 19702 29988 19740
rect 30156 19794 30212 19806
rect 30156 19742 30158 19794
rect 30210 19742 30212 19794
rect 29708 19618 29764 19628
rect 30156 19236 30212 19742
rect 31052 19794 31108 19806
rect 31052 19742 31054 19794
rect 31106 19742 31108 19794
rect 31052 19684 31108 19742
rect 30156 19170 30212 19180
rect 30268 19346 30324 19358
rect 30268 19294 30270 19346
rect 30322 19294 30324 19346
rect 29260 18958 29262 19010
rect 29314 18958 29316 19010
rect 29260 18900 29316 18958
rect 29036 18844 29316 18900
rect 28028 18174 28030 18226
rect 28082 18174 28084 18226
rect 28028 18162 28084 18174
rect 28252 18338 28308 18350
rect 28252 18286 28254 18338
rect 28306 18286 28308 18338
rect 28028 17890 28084 17902
rect 28028 17838 28030 17890
rect 28082 17838 28084 17890
rect 28028 17778 28084 17838
rect 28252 17890 28308 18286
rect 28252 17838 28254 17890
rect 28306 17838 28308 17890
rect 28252 17826 28308 17838
rect 28700 18338 28756 18350
rect 28700 18286 28702 18338
rect 28754 18286 28756 18338
rect 28028 17726 28030 17778
rect 28082 17726 28084 17778
rect 28028 17444 28084 17726
rect 28028 17378 28084 17388
rect 28476 17442 28532 17454
rect 28476 17390 28478 17442
rect 28530 17390 28532 17442
rect 28476 17332 28532 17390
rect 28476 17266 28532 17276
rect 27804 16930 27860 16940
rect 28476 16996 28532 17006
rect 27132 15934 27134 15986
rect 27186 15934 27188 15986
rect 26908 15876 26964 15886
rect 26908 15782 26964 15820
rect 26684 15262 26686 15314
rect 26738 15262 26740 15314
rect 26684 15250 26740 15262
rect 26908 15316 26964 15326
rect 26124 14802 26180 14812
rect 26236 14644 26292 14654
rect 26124 14532 26180 14542
rect 26124 14438 26180 14476
rect 25564 13916 25732 13972
rect 25340 13804 25620 13860
rect 24780 12962 24836 13020
rect 25452 13636 25508 13646
rect 24780 12910 24782 12962
rect 24834 12910 24836 12962
rect 24780 12898 24836 12910
rect 25228 12962 25284 12974
rect 25228 12910 25230 12962
rect 25282 12910 25284 12962
rect 25228 12852 25284 12910
rect 25228 12786 25284 12796
rect 25340 12964 25396 12974
rect 25228 12180 25284 12190
rect 25228 12086 25284 12124
rect 24556 12068 24612 12078
rect 24612 12012 24724 12068
rect 24556 12002 24612 12012
rect 24444 11190 24500 11228
rect 23772 10658 23828 10668
rect 24332 9828 24388 9838
rect 24332 9734 24388 9772
rect 24668 9268 24724 12012
rect 25340 11506 25396 12908
rect 25340 11454 25342 11506
rect 25394 11454 25396 11506
rect 25340 11442 25396 11454
rect 25452 12852 25508 13580
rect 25452 12180 25508 12796
rect 25452 11394 25508 12124
rect 25452 11342 25454 11394
rect 25506 11342 25508 11394
rect 25116 11282 25172 11294
rect 25116 11230 25118 11282
rect 25170 11230 25172 11282
rect 25004 10388 25060 10398
rect 24780 9940 24836 9950
rect 24780 9826 24836 9884
rect 24780 9774 24782 9826
rect 24834 9774 24836 9826
rect 24780 9762 24836 9774
rect 25004 9826 25060 10332
rect 25116 10052 25172 11230
rect 25228 11284 25284 11294
rect 25228 10610 25284 11228
rect 25340 10724 25396 10734
rect 25340 10630 25396 10668
rect 25228 10558 25230 10610
rect 25282 10558 25284 10610
rect 25228 10546 25284 10558
rect 25116 9986 25172 9996
rect 25004 9774 25006 9826
rect 25058 9774 25060 9826
rect 25004 9762 25060 9774
rect 25452 9828 25508 11342
rect 25452 9762 25508 9772
rect 24892 9602 24948 9614
rect 24892 9550 24894 9602
rect 24946 9550 24948 9602
rect 24780 9268 24836 9278
rect 24668 9212 24780 9268
rect 24780 9174 24836 9212
rect 24892 8148 24948 9550
rect 25228 9604 25284 9614
rect 25228 9510 25284 9548
rect 24444 8092 24948 8148
rect 25340 8818 25396 8830
rect 25340 8766 25342 8818
rect 25394 8766 25396 8818
rect 23436 7588 23492 7598
rect 23436 7494 23492 7532
rect 23772 7588 23828 7598
rect 23772 7494 23828 7532
rect 23772 6692 23828 6702
rect 23772 6598 23828 6636
rect 24444 6690 24500 8092
rect 25116 8036 25172 8046
rect 25116 7942 25172 7980
rect 25340 7588 25396 8766
rect 25340 7522 25396 7532
rect 25564 7250 25620 13804
rect 25676 13748 25732 13916
rect 25900 13748 25956 13758
rect 25676 13746 25956 13748
rect 25676 13694 25902 13746
rect 25954 13694 25956 13746
rect 25676 13692 25956 13694
rect 25676 13076 25732 13086
rect 25732 13020 25844 13076
rect 25676 13010 25732 13020
rect 25788 12290 25844 13020
rect 25900 12740 25956 13692
rect 26236 13746 26292 14588
rect 26796 14530 26852 14542
rect 26796 14478 26798 14530
rect 26850 14478 26852 14530
rect 26460 14418 26516 14430
rect 26460 14366 26462 14418
rect 26514 14366 26516 14418
rect 26236 13694 26238 13746
rect 26290 13694 26292 13746
rect 26012 13188 26068 13198
rect 26012 13094 26068 13132
rect 26236 13188 26292 13694
rect 26236 13122 26292 13132
rect 26348 14306 26404 14318
rect 26348 14254 26350 14306
rect 26402 14254 26404 14306
rect 26348 12964 26404 14254
rect 26348 12898 26404 12908
rect 26012 12740 26068 12750
rect 25900 12684 26012 12740
rect 26012 12674 26068 12684
rect 25788 12238 25790 12290
rect 25842 12238 25844 12290
rect 25788 12226 25844 12238
rect 26460 11956 26516 14366
rect 26572 14420 26628 14430
rect 26572 13970 26628 14364
rect 26572 13918 26574 13970
rect 26626 13918 26628 13970
rect 26572 13906 26628 13918
rect 26796 14308 26852 14478
rect 26908 14308 26964 15260
rect 27132 15148 27188 15934
rect 27244 15988 27300 15998
rect 27244 15894 27300 15932
rect 28140 15986 28196 15998
rect 28140 15934 28142 15986
rect 28194 15934 28196 15986
rect 27804 15876 27860 15886
rect 27356 15874 27860 15876
rect 27356 15822 27806 15874
rect 27858 15822 27860 15874
rect 27356 15820 27860 15822
rect 27244 15316 27300 15326
rect 27356 15316 27412 15820
rect 27804 15810 27860 15820
rect 28140 15876 28196 15934
rect 28140 15810 28196 15820
rect 28476 15428 28532 16940
rect 28700 16884 28756 18286
rect 28700 16790 28756 16828
rect 28812 18228 28868 18238
rect 29036 18228 29092 18844
rect 29148 18340 29204 18350
rect 29204 18284 29316 18340
rect 29148 18246 29204 18284
rect 28812 18226 29092 18228
rect 28812 18174 28814 18226
rect 28866 18174 29092 18226
rect 28812 18172 29092 18174
rect 28588 16100 28644 16110
rect 28588 16006 28644 16044
rect 27244 15314 27412 15316
rect 27244 15262 27246 15314
rect 27298 15262 27412 15314
rect 27244 15260 27412 15262
rect 28140 15372 28532 15428
rect 27244 15250 27300 15260
rect 27132 15092 27412 15148
rect 27132 14756 27188 14766
rect 27132 14642 27188 14700
rect 27132 14590 27134 14642
rect 27186 14590 27188 14642
rect 27132 14578 27188 14590
rect 27244 14644 27300 14654
rect 26796 14252 26964 14308
rect 26796 13972 26852 14252
rect 26908 13972 26964 14252
rect 27020 14532 27076 14542
rect 27020 14308 27076 14476
rect 27244 14530 27300 14588
rect 27244 14478 27246 14530
rect 27298 14478 27300 14530
rect 27244 14466 27300 14478
rect 27356 14530 27412 15092
rect 27580 14756 27636 14766
rect 27916 14756 27972 14766
rect 27636 14700 27860 14756
rect 27580 14690 27636 14700
rect 27804 14642 27860 14700
rect 27916 14662 27972 14700
rect 27804 14590 27806 14642
rect 27858 14590 27860 14642
rect 27804 14578 27860 14590
rect 28028 14644 28084 14654
rect 27356 14478 27358 14530
rect 27410 14478 27412 14530
rect 27356 14466 27412 14478
rect 27020 14214 27076 14252
rect 27916 14308 27972 14318
rect 27356 14196 27412 14206
rect 27412 14140 27524 14196
rect 27356 14130 27412 14140
rect 26908 13916 27412 13972
rect 26796 13906 26852 13916
rect 27356 13858 27412 13916
rect 27356 13806 27358 13858
rect 27410 13806 27412 13858
rect 27356 13794 27412 13806
rect 26796 13746 26852 13758
rect 26796 13694 26798 13746
rect 26850 13694 26852 13746
rect 26684 12962 26740 12974
rect 26684 12910 26686 12962
rect 26738 12910 26740 12962
rect 26684 12740 26740 12910
rect 26684 12068 26740 12684
rect 26684 12002 26740 12012
rect 26460 11890 26516 11900
rect 26796 10724 26852 13694
rect 27020 13746 27076 13758
rect 27020 13694 27022 13746
rect 27074 13694 27076 13746
rect 27020 13636 27076 13694
rect 27020 13412 27076 13580
rect 27020 13346 27076 13356
rect 27244 13746 27300 13758
rect 27244 13694 27246 13746
rect 27298 13694 27300 13746
rect 27244 13412 27300 13694
rect 27356 13636 27412 13646
rect 27468 13636 27524 14140
rect 27916 13972 27972 14252
rect 27804 13916 27972 13972
rect 27692 13748 27748 13758
rect 27356 13634 27524 13636
rect 27356 13582 27358 13634
rect 27410 13582 27524 13634
rect 27356 13580 27524 13582
rect 27580 13746 27748 13748
rect 27580 13694 27694 13746
rect 27746 13694 27748 13746
rect 27580 13692 27748 13694
rect 27356 13570 27412 13580
rect 27300 13356 27412 13412
rect 27244 13346 27300 13356
rect 26908 13188 26964 13198
rect 26908 13094 26964 13132
rect 27132 13076 27188 13086
rect 27132 12982 27188 13020
rect 27132 12740 27188 12750
rect 27020 12068 27076 12078
rect 27020 11974 27076 12012
rect 27132 11620 27188 12684
rect 27020 11564 27188 11620
rect 27244 11956 27300 11966
rect 27244 11618 27300 11900
rect 27244 11566 27246 11618
rect 27298 11566 27300 11618
rect 25676 10668 26852 10724
rect 26908 11508 26964 11518
rect 25676 9042 25732 10668
rect 25900 10498 25956 10510
rect 25900 10446 25902 10498
rect 25954 10446 25956 10498
rect 25900 10388 25956 10446
rect 26572 10388 26628 10398
rect 25900 10322 25956 10332
rect 26460 10386 26628 10388
rect 26460 10334 26574 10386
rect 26626 10334 26628 10386
rect 26460 10332 26628 10334
rect 26460 9940 26516 10332
rect 26572 10322 26628 10332
rect 26460 9874 26516 9884
rect 26572 9828 26628 9838
rect 26908 9828 26964 11452
rect 27020 10722 27076 11564
rect 27244 11554 27300 11566
rect 27356 11506 27412 13356
rect 27468 13076 27524 13086
rect 27468 12404 27524 13020
rect 27580 12852 27636 13692
rect 27692 13682 27748 13692
rect 27804 13524 27860 13916
rect 27580 12758 27636 12796
rect 27692 13468 27860 13524
rect 27916 13634 27972 13646
rect 27916 13582 27918 13634
rect 27970 13582 27972 13634
rect 27580 12404 27636 12414
rect 27468 12402 27636 12404
rect 27468 12350 27582 12402
rect 27634 12350 27636 12402
rect 27468 12348 27636 12350
rect 27580 12338 27636 12348
rect 27356 11454 27358 11506
rect 27410 11454 27412 11506
rect 27356 11442 27412 11454
rect 27692 11508 27748 13468
rect 27804 12964 27860 12974
rect 27804 12870 27860 12908
rect 27692 11414 27748 11452
rect 27804 11618 27860 11630
rect 27804 11566 27806 11618
rect 27858 11566 27860 11618
rect 27804 11172 27860 11566
rect 27916 11394 27972 13582
rect 28028 13636 28084 14588
rect 28140 14084 28196 15372
rect 28252 14420 28308 14430
rect 28252 14326 28308 14364
rect 28364 14308 28420 14318
rect 28588 14308 28644 14318
rect 28364 14214 28420 14252
rect 28476 14306 28644 14308
rect 28476 14254 28590 14306
rect 28642 14254 28644 14306
rect 28476 14252 28644 14254
rect 28140 14028 28420 14084
rect 28140 13860 28196 13870
rect 28140 13766 28196 13804
rect 28028 13570 28084 13580
rect 28252 13746 28308 13758
rect 28252 13694 28254 13746
rect 28306 13694 28308 13746
rect 28140 13412 28196 13422
rect 28252 13412 28308 13694
rect 28196 13356 28308 13412
rect 28140 13346 28196 13356
rect 28364 13300 28420 14028
rect 28252 13244 28420 13300
rect 28028 13188 28084 13198
rect 28028 12962 28084 13132
rect 28028 12910 28030 12962
rect 28082 12910 28084 12962
rect 28028 12898 28084 12910
rect 28140 12740 28196 12750
rect 28140 12646 28196 12684
rect 28252 12738 28308 13244
rect 28252 12686 28254 12738
rect 28306 12686 28308 12738
rect 27916 11342 27918 11394
rect 27970 11342 27972 11394
rect 27916 11330 27972 11342
rect 28028 12628 28084 12638
rect 27244 11116 27860 11172
rect 27020 10670 27022 10722
rect 27074 10670 27076 10722
rect 27020 10658 27076 10670
rect 27132 10724 27188 10734
rect 27244 10724 27300 11116
rect 27132 10722 27300 10724
rect 27132 10670 27134 10722
rect 27186 10670 27300 10722
rect 27132 10668 27300 10670
rect 27132 10658 27188 10668
rect 27356 10610 27412 10622
rect 27356 10558 27358 10610
rect 27410 10558 27412 10610
rect 27132 10052 27188 10062
rect 27020 9828 27076 9838
rect 26908 9772 27020 9828
rect 26572 9734 26628 9772
rect 26012 9716 26068 9726
rect 25676 8990 25678 9042
rect 25730 8990 25732 9042
rect 25676 8482 25732 8990
rect 25676 8430 25678 8482
rect 25730 8430 25732 8482
rect 25676 8418 25732 8430
rect 25900 9714 26068 9716
rect 25900 9662 26014 9714
rect 26066 9662 26068 9714
rect 25900 9660 26068 9662
rect 25900 9380 25956 9660
rect 26012 9650 26068 9660
rect 25900 8260 25956 9324
rect 26796 9604 26852 9614
rect 26012 9268 26068 9278
rect 26012 9154 26068 9212
rect 26796 9266 26852 9548
rect 26796 9214 26798 9266
rect 26850 9214 26852 9266
rect 26796 9202 26852 9214
rect 26012 9102 26014 9154
rect 26066 9102 26068 9154
rect 26012 9090 26068 9102
rect 26460 9156 26516 9166
rect 26460 9062 26516 9100
rect 26908 9156 26964 9166
rect 25564 7198 25566 7250
rect 25618 7198 25620 7250
rect 25564 7186 25620 7198
rect 25676 8204 25956 8260
rect 26348 8258 26404 8270
rect 26348 8206 26350 8258
rect 26402 8206 26404 8258
rect 24444 6638 24446 6690
rect 24498 6638 24500 6690
rect 24444 6626 24500 6638
rect 25676 3666 25732 8204
rect 26012 8146 26068 8158
rect 26012 8094 26014 8146
rect 26066 8094 26068 8146
rect 25900 8036 25956 8046
rect 25900 7942 25956 7980
rect 26012 7700 26068 8094
rect 26236 7700 26292 7710
rect 26348 7700 26404 8206
rect 26012 7698 26404 7700
rect 26012 7646 26238 7698
rect 26290 7646 26404 7698
rect 26012 7644 26404 7646
rect 26908 7698 26964 9100
rect 26908 7646 26910 7698
rect 26962 7646 26964 7698
rect 25788 7362 25844 7374
rect 25788 7310 25790 7362
rect 25842 7310 25844 7362
rect 25788 6692 25844 7310
rect 25788 6626 25844 6636
rect 26012 6468 26068 7644
rect 26236 7634 26292 7644
rect 26908 7634 26964 7646
rect 27020 9154 27076 9772
rect 27020 9102 27022 9154
rect 27074 9102 27076 9154
rect 26012 6402 26068 6412
rect 26460 7250 26516 7262
rect 26460 7198 26462 7250
rect 26514 7198 26516 7250
rect 26348 4228 26404 4238
rect 25676 3614 25678 3666
rect 25730 3614 25732 3666
rect 25676 3602 25732 3614
rect 26124 4226 26404 4228
rect 26124 4174 26350 4226
rect 26402 4174 26404 4226
rect 26124 4172 26404 4174
rect 23548 3556 23604 3566
rect 23548 3462 23604 3500
rect 26124 3554 26180 4172
rect 26348 4162 26404 4172
rect 26124 3502 26126 3554
rect 26178 3502 26180 3554
rect 23324 3390 23326 3442
rect 23378 3390 23380 3442
rect 23324 3378 23380 3390
rect 26124 3388 26180 3502
rect 26460 3554 26516 7198
rect 27020 6916 27076 9102
rect 27132 9492 27188 9996
rect 27132 9154 27188 9436
rect 27356 9266 27412 10558
rect 28028 10610 28084 12572
rect 28252 11956 28308 12686
rect 28140 11900 28308 11956
rect 28364 12964 28420 12974
rect 28140 11172 28196 11900
rect 28252 11732 28308 11742
rect 28252 11618 28308 11676
rect 28252 11566 28254 11618
rect 28306 11566 28308 11618
rect 28252 11554 28308 11566
rect 28252 11172 28308 11182
rect 28140 11116 28252 11172
rect 28252 11106 28308 11116
rect 28140 10724 28196 10734
rect 28364 10724 28420 12908
rect 28476 12180 28532 14252
rect 28588 14242 28644 14252
rect 28812 12628 28868 18172
rect 29260 17668 29316 18284
rect 29708 18338 29764 18350
rect 29708 18286 29710 18338
rect 29762 18286 29764 18338
rect 29708 17892 29764 18286
rect 30044 18338 30100 18350
rect 30044 18286 30046 18338
rect 30098 18286 30100 18338
rect 29708 17836 29988 17892
rect 29372 17780 29428 17790
rect 29372 17686 29428 17724
rect 29260 16770 29316 17612
rect 29708 17668 29764 17678
rect 29708 17574 29764 17612
rect 29260 16718 29262 16770
rect 29314 16718 29316 16770
rect 29260 16100 29316 16718
rect 29260 16034 29316 16044
rect 29484 17442 29540 17454
rect 29484 17390 29486 17442
rect 29538 17390 29540 17442
rect 29260 15876 29316 15886
rect 29260 15782 29316 15820
rect 29484 15538 29540 17390
rect 29820 17332 29876 17342
rect 29820 16996 29876 17276
rect 29596 16100 29652 16110
rect 29596 16006 29652 16044
rect 29820 15986 29876 16940
rect 29820 15934 29822 15986
rect 29874 15934 29876 15986
rect 29820 15652 29876 15934
rect 29932 15988 29988 17836
rect 30044 17780 30100 18286
rect 30044 17714 30100 17724
rect 30268 18228 30324 19294
rect 30716 19236 30772 19246
rect 30716 19142 30772 19180
rect 31052 19124 31108 19628
rect 31164 19346 31220 20750
rect 31276 20580 31332 22316
rect 31500 21812 31556 21822
rect 31500 21026 31556 21756
rect 31836 21588 31892 23324
rect 31948 21700 32004 25676
rect 32172 25508 32228 26238
rect 32060 25452 32228 25508
rect 32060 25282 32116 25452
rect 32060 25230 32062 25282
rect 32114 25230 32116 25282
rect 32060 24500 32116 25230
rect 32172 25282 32228 25294
rect 32172 25230 32174 25282
rect 32226 25230 32228 25282
rect 32172 24722 32228 25230
rect 32284 25284 32340 25294
rect 32396 25284 32452 26684
rect 32508 26516 32564 26526
rect 32508 26402 32564 26460
rect 32508 26350 32510 26402
rect 32562 26350 32564 26402
rect 32508 26338 32564 26350
rect 32956 26290 33012 26302
rect 32956 26238 32958 26290
rect 33010 26238 33012 26290
rect 32844 26180 32900 26190
rect 32732 26124 32844 26180
rect 32284 25282 32452 25284
rect 32284 25230 32286 25282
rect 32338 25230 32452 25282
rect 32284 25228 32452 25230
rect 32284 25218 32340 25228
rect 32172 24670 32174 24722
rect 32226 24670 32228 24722
rect 32172 24658 32228 24670
rect 32060 24434 32116 24444
rect 32396 23940 32452 25228
rect 32508 25284 32564 25294
rect 32508 25190 32564 25228
rect 32172 23380 32228 23390
rect 32172 23154 32228 23324
rect 32172 23102 32174 23154
rect 32226 23102 32228 23154
rect 32172 23090 32228 23102
rect 32284 22260 32340 22270
rect 32284 22166 32340 22204
rect 32396 22036 32452 23884
rect 32284 21980 32452 22036
rect 32172 21700 32228 21710
rect 31948 21698 32228 21700
rect 31948 21646 32174 21698
rect 32226 21646 32228 21698
rect 31948 21644 32228 21646
rect 31836 21532 32004 21588
rect 31500 20974 31502 21026
rect 31554 20974 31556 21026
rect 31500 20962 31556 20974
rect 31724 21474 31780 21486
rect 31724 21422 31726 21474
rect 31778 21422 31780 21474
rect 31724 20916 31780 21422
rect 31836 21364 31892 21374
rect 31836 21270 31892 21308
rect 31948 21140 32004 21532
rect 31724 20850 31780 20860
rect 31836 21084 32004 21140
rect 31276 20514 31332 20524
rect 31500 20020 31556 20030
rect 31500 19906 31556 19964
rect 31500 19854 31502 19906
rect 31554 19854 31556 19906
rect 31164 19294 31166 19346
rect 31218 19294 31220 19346
rect 31164 19282 31220 19294
rect 31276 19796 31332 19806
rect 31052 19030 31108 19068
rect 31276 19012 31332 19740
rect 31276 19010 31444 19012
rect 31276 18958 31278 19010
rect 31330 18958 31444 19010
rect 31276 18956 31444 18958
rect 31276 18946 31332 18956
rect 31164 18900 31220 18910
rect 30716 18340 30772 18350
rect 31164 18340 31220 18844
rect 30716 18338 31220 18340
rect 30716 18286 30718 18338
rect 30770 18286 31166 18338
rect 31218 18286 31220 18338
rect 30716 18284 31220 18286
rect 31388 18340 31444 18956
rect 31500 19010 31556 19854
rect 31500 18958 31502 19010
rect 31554 18958 31556 19010
rect 31500 18900 31556 18958
rect 31500 18834 31556 18844
rect 31724 18340 31780 18350
rect 31388 18284 31724 18340
rect 30716 18228 30772 18284
rect 31164 18274 31220 18284
rect 31724 18246 31780 18284
rect 30268 18172 30772 18228
rect 31276 18226 31332 18238
rect 31276 18174 31278 18226
rect 31330 18174 31332 18226
rect 30268 17444 30324 18172
rect 30380 17668 30436 17678
rect 30380 17666 31220 17668
rect 30380 17614 30382 17666
rect 30434 17614 31220 17666
rect 30380 17612 31220 17614
rect 30380 17602 30436 17612
rect 30268 17388 30436 17444
rect 29932 15922 29988 15932
rect 30268 16100 30324 16110
rect 29820 15586 29876 15596
rect 29484 15486 29486 15538
rect 29538 15486 29540 15538
rect 29484 15474 29540 15486
rect 30268 15540 30324 16044
rect 30380 15988 30436 17388
rect 31164 16210 31220 17612
rect 31164 16158 31166 16210
rect 31218 16158 31220 16210
rect 31164 16146 31220 16158
rect 31276 16098 31332 18174
rect 31276 16046 31278 16098
rect 31330 16046 31332 16098
rect 31276 16034 31332 16046
rect 31388 17668 31444 17678
rect 31388 16884 31444 17612
rect 31052 15988 31108 15998
rect 30380 15986 30660 15988
rect 30380 15934 30382 15986
rect 30434 15934 30660 15986
rect 30380 15932 30660 15934
rect 30380 15922 30436 15932
rect 30268 15538 30548 15540
rect 30268 15486 30270 15538
rect 30322 15486 30548 15538
rect 30268 15484 30548 15486
rect 30268 15474 30324 15484
rect 30492 15426 30548 15484
rect 30492 15374 30494 15426
rect 30546 15374 30548 15426
rect 30492 15362 30548 15374
rect 30604 14868 30660 15932
rect 31108 15932 31220 15988
rect 31052 15894 31108 15932
rect 30604 14802 30660 14812
rect 30716 15876 30772 15886
rect 30716 15538 30772 15820
rect 30716 15486 30718 15538
rect 30770 15486 30772 15538
rect 30716 14644 30772 15486
rect 31164 15428 31220 15932
rect 31164 15362 31220 15372
rect 30940 15314 30996 15326
rect 30940 15262 30942 15314
rect 30994 15262 30996 15314
rect 30828 15204 30884 15242
rect 30828 15138 30884 15148
rect 30940 14756 30996 15262
rect 31052 15316 31108 15326
rect 31052 15222 31108 15260
rect 30044 14588 30660 14644
rect 29708 14532 29764 14542
rect 29708 14438 29764 14476
rect 30044 14530 30100 14588
rect 30044 14478 30046 14530
rect 30098 14478 30100 14530
rect 30044 14466 30100 14478
rect 30604 14530 30660 14588
rect 30716 14578 30772 14588
rect 30828 14700 30996 14756
rect 31052 15092 31108 15102
rect 30604 14478 30606 14530
rect 30658 14478 30660 14530
rect 28924 14420 28980 14430
rect 28924 13746 28980 14364
rect 30156 14418 30212 14430
rect 30492 14420 30548 14430
rect 30156 14366 30158 14418
rect 30210 14366 30212 14418
rect 28924 13694 28926 13746
rect 28978 13694 28980 13746
rect 28924 13682 28980 13694
rect 29148 13860 29204 13870
rect 30044 13860 30100 13870
rect 29148 12964 29204 13804
rect 29484 13858 30100 13860
rect 29484 13806 30046 13858
rect 30098 13806 30100 13858
rect 29484 13804 30100 13806
rect 29484 13300 29540 13804
rect 30044 13794 30100 13804
rect 29260 13244 29540 13300
rect 29596 13412 29652 13422
rect 30156 13412 30212 14366
rect 30268 14418 30548 14420
rect 30268 14366 30494 14418
rect 30546 14366 30548 14418
rect 30268 14364 30548 14366
rect 30268 13746 30324 14364
rect 30492 14354 30548 14364
rect 30268 13694 30270 13746
rect 30322 13694 30324 13746
rect 30268 13682 30324 13694
rect 30604 13860 30660 14478
rect 30380 13524 30436 13534
rect 30156 13356 30324 13412
rect 29260 13074 29316 13244
rect 29260 13022 29262 13074
rect 29314 13022 29316 13074
rect 29260 13010 29316 13022
rect 28812 12562 28868 12572
rect 28924 12962 29204 12964
rect 28924 12910 29150 12962
rect 29202 12910 29204 12962
rect 28924 12908 29204 12910
rect 28924 12292 28980 12908
rect 29148 12898 29204 12908
rect 29372 12738 29428 12750
rect 29372 12686 29374 12738
rect 29426 12686 29428 12738
rect 29372 12628 29428 12686
rect 29372 12562 29428 12572
rect 29596 12404 29652 13356
rect 28924 12198 28980 12236
rect 29484 12348 29652 12404
rect 29708 13188 29764 13198
rect 30156 13188 30212 13198
rect 29484 12180 29540 12348
rect 28476 12086 28532 12124
rect 29148 12178 29540 12180
rect 29148 12126 29486 12178
rect 29538 12126 29540 12178
rect 29148 12124 29540 12126
rect 28812 12066 28868 12078
rect 28812 12014 28814 12066
rect 28866 12014 28868 12066
rect 28476 11396 28532 11406
rect 28476 11302 28532 11340
rect 28140 10722 28364 10724
rect 28140 10670 28142 10722
rect 28194 10670 28364 10722
rect 28140 10668 28364 10670
rect 28140 10658 28196 10668
rect 28364 10630 28420 10668
rect 28812 10722 28868 12014
rect 28812 10670 28814 10722
rect 28866 10670 28868 10722
rect 28812 10658 28868 10670
rect 28028 10558 28030 10610
rect 28082 10558 28084 10610
rect 27356 9214 27358 9266
rect 27410 9214 27412 9266
rect 27356 9202 27412 9214
rect 27580 10052 27636 10062
rect 27580 9266 27636 9996
rect 28028 9828 28084 10558
rect 28924 10610 28980 10622
rect 28924 10558 28926 10610
rect 28978 10558 28980 10610
rect 27692 9772 27972 9828
rect 28028 9772 28532 9828
rect 27692 9714 27748 9772
rect 27692 9662 27694 9714
rect 27746 9662 27748 9714
rect 27692 9650 27748 9662
rect 27580 9214 27582 9266
rect 27634 9214 27636 9266
rect 27580 9202 27636 9214
rect 27804 9602 27860 9614
rect 27804 9550 27806 9602
rect 27858 9550 27860 9602
rect 27132 9102 27134 9154
rect 27186 9102 27188 9154
rect 27132 9090 27188 9102
rect 27692 9156 27748 9166
rect 27804 9156 27860 9550
rect 27692 9154 27860 9156
rect 27692 9102 27694 9154
rect 27746 9102 27860 9154
rect 27692 9100 27860 9102
rect 27692 9090 27748 9100
rect 27916 8596 27972 9772
rect 28476 9714 28532 9772
rect 28476 9662 28478 9714
rect 28530 9662 28532 9714
rect 28252 9602 28308 9614
rect 28252 9550 28254 9602
rect 28306 9550 28308 9602
rect 28252 8708 28308 9550
rect 28476 9156 28532 9662
rect 28588 9716 28644 9726
rect 28588 9714 28756 9716
rect 28588 9662 28590 9714
rect 28642 9662 28756 9714
rect 28588 9660 28756 9662
rect 28588 9650 28644 9660
rect 28588 9156 28644 9166
rect 28532 9154 28644 9156
rect 28532 9102 28590 9154
rect 28642 9102 28644 9154
rect 28532 9100 28644 9102
rect 28476 9062 28532 9100
rect 28588 9090 28644 9100
rect 28700 9044 28756 9660
rect 28924 9268 28980 10558
rect 28924 9202 28980 9212
rect 29148 10050 29204 12124
rect 29484 12114 29540 12124
rect 29596 12180 29652 12190
rect 29484 11732 29540 11742
rect 29148 9998 29150 10050
rect 29202 9998 29204 10050
rect 29148 9044 29204 9998
rect 29260 11172 29316 11182
rect 29484 11172 29540 11676
rect 29596 11394 29652 12124
rect 29708 11506 29764 13132
rect 29820 13186 30212 13188
rect 29820 13134 30158 13186
rect 30210 13134 30212 13186
rect 29820 13132 30212 13134
rect 29820 12962 29876 13132
rect 30156 13122 30212 13132
rect 29820 12910 29822 12962
rect 29874 12910 29876 12962
rect 29820 12898 29876 12910
rect 30044 12964 30100 12974
rect 30268 12964 30324 13356
rect 30044 12962 30324 12964
rect 30044 12910 30046 12962
rect 30098 12910 30324 12962
rect 30044 12908 30324 12910
rect 30044 12898 30100 12908
rect 30380 12852 30436 13468
rect 30156 12796 30436 12852
rect 30492 13188 30548 13198
rect 30156 12738 30212 12796
rect 30492 12740 30548 13132
rect 30156 12686 30158 12738
rect 30210 12686 30212 12738
rect 29708 11454 29710 11506
rect 29762 11454 29764 11506
rect 29708 11442 29764 11454
rect 29932 12292 29988 12302
rect 29596 11342 29598 11394
rect 29650 11342 29652 11394
rect 29596 11330 29652 11342
rect 29820 11396 29876 11406
rect 29484 11116 29764 11172
rect 29260 9828 29316 11116
rect 29708 10050 29764 11116
rect 29708 9998 29710 10050
rect 29762 9998 29764 10050
rect 29708 9986 29764 9998
rect 29820 10052 29876 11340
rect 29932 11394 29988 12236
rect 29932 11342 29934 11394
rect 29986 11342 29988 11394
rect 29932 11330 29988 11342
rect 30044 12180 30100 12190
rect 30044 11394 30100 12124
rect 30044 11342 30046 11394
rect 30098 11342 30100 11394
rect 30044 11330 30100 11342
rect 30156 11172 30212 12686
rect 30380 12684 30548 12740
rect 30380 11956 30436 12684
rect 30604 12628 30660 13804
rect 30716 13858 30772 13870
rect 30716 13806 30718 13858
rect 30770 13806 30772 13858
rect 30716 13076 30772 13806
rect 30828 13188 30884 14700
rect 30940 14530 30996 14542
rect 30940 14478 30942 14530
rect 30994 14478 30996 14530
rect 30940 14308 30996 14478
rect 30940 13748 30996 14252
rect 30940 13682 30996 13692
rect 31052 14532 31108 15036
rect 31052 13746 31108 14476
rect 31052 13694 31054 13746
rect 31106 13694 31108 13746
rect 31052 13682 31108 13694
rect 31164 13634 31220 13646
rect 31164 13582 31166 13634
rect 31218 13582 31220 13634
rect 31164 13524 31220 13582
rect 31164 13458 31220 13468
rect 30828 13122 30884 13132
rect 31276 13186 31332 13198
rect 31276 13134 31278 13186
rect 31330 13134 31332 13186
rect 30716 13010 30772 13020
rect 30828 12852 30884 12862
rect 30492 12572 30604 12628
rect 30492 12178 30548 12572
rect 30604 12562 30660 12572
rect 30716 12850 30884 12852
rect 30716 12798 30830 12850
rect 30882 12798 30884 12850
rect 30716 12796 30884 12798
rect 30716 12402 30772 12796
rect 30828 12786 30884 12796
rect 30716 12350 30718 12402
rect 30770 12350 30772 12402
rect 30492 12126 30494 12178
rect 30546 12126 30548 12178
rect 30492 12114 30548 12126
rect 30604 12292 30660 12302
rect 30604 11956 30660 12236
rect 30716 12180 30772 12350
rect 30716 12114 30772 12124
rect 30940 12738 30996 12750
rect 31164 12740 31220 12750
rect 30940 12686 30942 12738
rect 30994 12686 30996 12738
rect 30380 11900 30660 11956
rect 30828 12068 30884 12078
rect 30828 11620 30884 12012
rect 30492 11564 30884 11620
rect 29932 11116 30212 11172
rect 30380 11396 30436 11406
rect 29932 10612 29988 11116
rect 30044 10836 30100 10846
rect 30044 10834 30212 10836
rect 30044 10782 30046 10834
rect 30098 10782 30212 10834
rect 30044 10780 30212 10782
rect 30044 10770 30100 10780
rect 29932 10610 30100 10612
rect 29932 10558 29934 10610
rect 29986 10558 30100 10610
rect 29932 10556 30100 10558
rect 29932 10546 29988 10556
rect 29932 10052 29988 10062
rect 29820 10050 29988 10052
rect 29820 9998 29934 10050
rect 29986 9998 29988 10050
rect 29820 9996 29988 9998
rect 29932 9986 29988 9996
rect 30044 10052 30100 10556
rect 30156 10052 30212 10780
rect 30380 10834 30436 11340
rect 30492 11394 30548 11564
rect 30940 11508 30996 12686
rect 30492 11342 30494 11394
rect 30546 11342 30548 11394
rect 30492 11330 30548 11342
rect 30716 11452 30940 11508
rect 30380 10782 30382 10834
rect 30434 10782 30436 10834
rect 30380 10770 30436 10782
rect 30604 11284 30660 11294
rect 30492 10724 30548 10734
rect 30604 10724 30660 11228
rect 30492 10722 30660 10724
rect 30492 10670 30494 10722
rect 30546 10670 30660 10722
rect 30492 10668 30660 10670
rect 30492 10658 30548 10668
rect 30604 10388 30660 10398
rect 30156 9996 30436 10052
rect 30044 9986 30100 9996
rect 29260 9380 29316 9772
rect 30156 9828 30212 9838
rect 29372 9714 29428 9726
rect 29372 9662 29374 9714
rect 29426 9662 29428 9714
rect 29372 9492 29428 9662
rect 30044 9604 30100 9614
rect 30044 9510 30100 9548
rect 29372 9380 29428 9436
rect 29596 9380 29652 9390
rect 29372 9324 29596 9380
rect 29260 9314 29316 9324
rect 29596 9314 29652 9324
rect 28700 9042 29204 9044
rect 28700 8990 29150 9042
rect 29202 8990 29204 9042
rect 28700 8988 29204 8990
rect 28252 8652 28532 8708
rect 27916 8540 28308 8596
rect 28140 8260 28196 8270
rect 27468 8148 27524 8158
rect 27468 7698 27524 8092
rect 28028 8148 28084 8158
rect 28028 8054 28084 8092
rect 27916 8036 27972 8046
rect 27468 7646 27470 7698
rect 27522 7646 27524 7698
rect 27468 7634 27524 7646
rect 27804 8034 27972 8036
rect 27804 7982 27918 8034
rect 27970 7982 27972 8034
rect 27804 7980 27972 7982
rect 27468 6916 27524 6926
rect 27020 6914 27524 6916
rect 27020 6862 27470 6914
rect 27522 6862 27524 6914
rect 27020 6860 27524 6862
rect 27468 6850 27524 6860
rect 26796 6580 26852 6590
rect 26796 6466 26852 6524
rect 27804 6580 27860 7980
rect 27916 7970 27972 7980
rect 27916 7700 27972 7710
rect 28140 7700 28196 8204
rect 28252 8258 28308 8540
rect 28252 8206 28254 8258
rect 28306 8206 28308 8258
rect 28252 8194 28308 8206
rect 28476 8146 28532 8652
rect 29148 8260 29204 8988
rect 29148 8194 29204 8204
rect 29372 9156 29428 9166
rect 29372 8372 29428 9100
rect 29372 8258 29428 8316
rect 29372 8206 29374 8258
rect 29426 8206 29428 8258
rect 29372 8194 29428 8206
rect 29708 8820 29764 8830
rect 29708 8258 29764 8764
rect 30156 8370 30212 9772
rect 30380 9826 30436 9996
rect 30380 9774 30382 9826
rect 30434 9774 30436 9826
rect 30380 9762 30436 9774
rect 30604 9826 30660 10332
rect 30604 9774 30606 9826
rect 30658 9774 30660 9826
rect 30604 9762 30660 9774
rect 30716 9716 30772 11452
rect 30940 11442 30996 11452
rect 31052 12738 31220 12740
rect 31052 12686 31166 12738
rect 31218 12686 31220 12738
rect 31052 12684 31220 12686
rect 30940 11282 30996 11294
rect 30940 11230 30942 11282
rect 30994 11230 30996 11282
rect 30940 10836 30996 11230
rect 31052 11284 31108 12684
rect 31164 12674 31220 12684
rect 31276 12290 31332 13134
rect 31276 12238 31278 12290
rect 31330 12238 31332 12290
rect 31276 12226 31332 12238
rect 31388 13076 31444 16828
rect 31724 16660 31780 16670
rect 31612 16100 31668 16110
rect 31612 15538 31668 16044
rect 31724 16098 31780 16604
rect 31724 16046 31726 16098
rect 31778 16046 31780 16098
rect 31724 16034 31780 16046
rect 31612 15486 31614 15538
rect 31666 15486 31668 15538
rect 31612 15474 31668 15486
rect 31500 15204 31556 15242
rect 31836 15148 31892 21084
rect 31948 20916 32004 20926
rect 32060 20916 32116 21644
rect 32172 21634 32228 21644
rect 31948 20914 32116 20916
rect 31948 20862 31950 20914
rect 32002 20862 32116 20914
rect 31948 20860 32116 20862
rect 31948 20850 32004 20860
rect 32060 20580 32116 20590
rect 31948 20020 32004 20030
rect 31948 19926 32004 19964
rect 32060 19010 32116 20524
rect 32284 20020 32340 21980
rect 32732 21812 32788 26124
rect 32844 26114 32900 26124
rect 32956 25732 33012 26238
rect 33180 26180 33236 27804
rect 33516 27300 33572 28590
rect 34300 28644 34356 28654
rect 34300 28550 34356 28588
rect 34636 28532 34692 29262
rect 34748 29092 34804 29374
rect 34748 29026 34804 29036
rect 34860 28868 34916 30940
rect 34972 30098 35028 33180
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 39564 31668 39620 31678
rect 39564 31574 39620 31612
rect 40012 31668 40068 31678
rect 39228 31554 39284 31566
rect 39228 31502 39230 31554
rect 39282 31502 39284 31554
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34972 30046 34974 30098
rect 35026 30046 35028 30098
rect 34972 30034 35028 30046
rect 35420 30436 35476 30446
rect 35196 29428 35252 29438
rect 35196 29334 35252 29372
rect 35420 29426 35476 30380
rect 35644 30324 35700 30334
rect 35644 30210 35700 30268
rect 39228 30324 39284 31502
rect 39900 31554 39956 31566
rect 39900 31502 39902 31554
rect 39954 31502 39956 31554
rect 39900 31444 39956 31502
rect 39900 31378 39956 31388
rect 39900 31220 39956 31230
rect 40012 31220 40068 31612
rect 39900 31218 40068 31220
rect 39900 31166 39902 31218
rect 39954 31166 40068 31218
rect 39900 31164 40068 31166
rect 40236 31554 40292 31566
rect 40236 31502 40238 31554
rect 40290 31502 40292 31554
rect 39900 31154 39956 31164
rect 40236 30996 40292 31502
rect 40236 30902 40292 30940
rect 39228 30258 39284 30268
rect 35644 30158 35646 30210
rect 35698 30158 35700 30210
rect 35644 30146 35700 30158
rect 35420 29374 35422 29426
rect 35474 29374 35476 29426
rect 35420 29362 35476 29374
rect 37100 29652 37156 29662
rect 34972 29316 35028 29326
rect 34972 29222 35028 29260
rect 35868 29316 35924 29326
rect 35868 29222 35924 29260
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 34748 28812 34916 28868
rect 35532 28868 35588 28878
rect 34748 28642 34804 28812
rect 34748 28590 34750 28642
rect 34802 28590 34804 28642
rect 34748 28578 34804 28590
rect 35420 28756 35476 28766
rect 35420 28642 35476 28700
rect 35532 28754 35588 28812
rect 35532 28702 35534 28754
rect 35586 28702 35588 28754
rect 35532 28690 35588 28702
rect 35420 28590 35422 28642
rect 35474 28590 35476 28642
rect 35420 28578 35476 28590
rect 36316 28644 36372 28654
rect 36316 28550 36372 28588
rect 37100 28644 37156 29596
rect 37100 28550 37156 28588
rect 37436 29428 37492 29438
rect 37436 28756 37492 29372
rect 39004 29428 39060 29438
rect 39004 29334 39060 29372
rect 40124 29314 40180 29326
rect 40124 29262 40126 29314
rect 40178 29262 40180 29314
rect 34636 28466 34692 28476
rect 34412 28420 34468 28430
rect 33740 27860 33796 27870
rect 33796 27804 33908 27860
rect 33740 27766 33796 27804
rect 33516 27234 33572 27244
rect 33852 27298 33908 27804
rect 34412 27858 34468 28364
rect 36092 28420 36148 28430
rect 36092 28326 36148 28364
rect 36988 28418 37044 28430
rect 36988 28366 36990 28418
rect 37042 28366 37044 28418
rect 36876 28084 36932 28094
rect 36988 28084 37044 28366
rect 36876 28082 37044 28084
rect 36876 28030 36878 28082
rect 36930 28030 37044 28082
rect 36876 28028 37044 28030
rect 37436 28082 37492 28700
rect 39900 29204 39956 29214
rect 37548 28644 37604 28654
rect 37548 28550 37604 28588
rect 39676 28642 39732 28654
rect 39676 28590 39678 28642
rect 39730 28590 39732 28642
rect 39676 28308 39732 28590
rect 39900 28530 39956 29148
rect 40124 28980 40180 29262
rect 40124 28914 40180 28924
rect 39900 28478 39902 28530
rect 39954 28478 39956 28530
rect 39900 28466 39956 28478
rect 40236 28642 40292 28654
rect 40236 28590 40238 28642
rect 40290 28590 40292 28642
rect 39676 28242 39732 28252
rect 40236 28308 40292 28590
rect 40236 28242 40292 28252
rect 37436 28030 37438 28082
rect 37490 28030 37492 28082
rect 36876 28018 36932 28028
rect 37436 28018 37492 28030
rect 34412 27806 34414 27858
rect 34466 27806 34468 27858
rect 34412 27794 34468 27806
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 33852 27246 33854 27298
rect 33906 27246 33908 27298
rect 33404 27188 33460 27198
rect 33404 27094 33460 27132
rect 33852 27186 33908 27246
rect 33852 27134 33854 27186
rect 33906 27134 33908 27186
rect 33852 27122 33908 27134
rect 34748 27300 34804 27310
rect 34748 27186 34804 27244
rect 34748 27134 34750 27186
rect 34802 27134 34804 27186
rect 34748 27122 34804 27134
rect 35196 27298 35252 27310
rect 35196 27246 35198 27298
rect 35250 27246 35252 27298
rect 35196 27186 35252 27246
rect 35196 27134 35198 27186
rect 35250 27134 35252 27186
rect 35196 27122 35252 27134
rect 34300 26850 34356 26862
rect 34300 26798 34302 26850
rect 34354 26798 34356 26850
rect 33404 26516 33460 26526
rect 33404 26422 33460 26460
rect 32956 25666 33012 25676
rect 33068 26124 33236 26180
rect 33292 26290 33348 26302
rect 33292 26238 33294 26290
rect 33346 26238 33348 26290
rect 33292 26180 33348 26238
rect 33964 26292 34020 26302
rect 34300 26292 34356 26798
rect 34412 26740 34468 26750
rect 34412 26514 34468 26684
rect 34412 26462 34414 26514
rect 34466 26462 34468 26514
rect 34412 26450 34468 26462
rect 34020 26236 34356 26292
rect 36540 26292 36596 26302
rect 33964 26198 34020 26236
rect 32844 25508 32900 25518
rect 33068 25508 33124 26124
rect 33292 26114 33348 26124
rect 33740 26180 33796 26190
rect 33740 26178 33908 26180
rect 33740 26126 33742 26178
rect 33794 26126 33908 26178
rect 33740 26124 33908 26126
rect 33740 26114 33796 26124
rect 33516 26068 33572 26078
rect 33292 25844 33348 25854
rect 33348 25788 33460 25844
rect 33292 25778 33348 25788
rect 32844 25506 33124 25508
rect 32844 25454 32846 25506
rect 32898 25454 33124 25506
rect 32844 25452 33124 25454
rect 33404 25506 33460 25788
rect 33404 25454 33406 25506
rect 33458 25454 33460 25506
rect 32844 22484 32900 25452
rect 33404 25442 33460 25454
rect 33516 25060 33572 26012
rect 33404 25004 33572 25060
rect 33068 24836 33124 24846
rect 33068 24742 33124 24780
rect 33180 24834 33236 24846
rect 33180 24782 33182 24834
rect 33234 24782 33236 24834
rect 33180 24724 33236 24782
rect 33180 24658 33236 24668
rect 33180 24498 33236 24510
rect 33180 24446 33182 24498
rect 33234 24446 33236 24498
rect 33068 23940 33124 23950
rect 33068 23846 33124 23884
rect 33180 23154 33236 24446
rect 33404 23716 33460 25004
rect 33852 24948 33908 26124
rect 33852 24892 34020 24948
rect 33516 24500 33572 24510
rect 33516 23938 33572 24444
rect 33964 24050 34020 24892
rect 33964 23998 33966 24050
rect 34018 23998 34020 24050
rect 33964 23986 34020 23998
rect 33516 23886 33518 23938
rect 33570 23886 33572 23938
rect 33516 23874 33572 23886
rect 33404 23660 33572 23716
rect 33292 23380 33348 23390
rect 33292 23286 33348 23324
rect 33180 23102 33182 23154
rect 33234 23102 33236 23154
rect 33180 23090 33236 23102
rect 32844 22418 32900 22428
rect 32956 22372 33012 22382
rect 32956 22278 33012 22316
rect 33180 22370 33236 22382
rect 33180 22318 33182 22370
rect 33234 22318 33236 22370
rect 33180 22036 33236 22318
rect 33516 22372 33572 23660
rect 34076 23604 34132 26236
rect 34860 26178 34916 26190
rect 34860 26126 34862 26178
rect 34914 26126 34916 26178
rect 34860 25732 34916 26126
rect 35308 26178 35364 26190
rect 35308 26126 35310 26178
rect 35362 26126 35364 26178
rect 35308 26068 35364 26126
rect 35308 26002 35364 26012
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35756 25732 35812 25742
rect 34860 25666 34916 25676
rect 35644 25676 35756 25732
rect 34636 24836 34692 24846
rect 34188 24724 34244 24734
rect 34188 24498 34244 24668
rect 34188 24446 34190 24498
rect 34242 24446 34244 24498
rect 34188 23938 34244 24446
rect 34188 23886 34190 23938
rect 34242 23886 34244 23938
rect 34188 23874 34244 23886
rect 34300 24722 34356 24734
rect 34300 24670 34302 24722
rect 34354 24670 34356 24722
rect 34300 23940 34356 24670
rect 34412 24612 34468 24622
rect 34412 24518 34468 24556
rect 34300 23874 34356 23884
rect 34636 23940 34692 24780
rect 35644 24722 35700 25676
rect 35756 25666 35812 25676
rect 36540 25732 36596 26236
rect 39004 26292 39060 26302
rect 39004 26198 39060 26236
rect 36540 25638 36596 25676
rect 40124 26178 40180 26190
rect 40124 26126 40126 26178
rect 40178 26126 40180 26178
rect 40124 25620 40180 26126
rect 40124 25554 40180 25564
rect 39004 25508 39060 25518
rect 39004 25414 39060 25452
rect 35756 25284 35812 25294
rect 35980 25284 36036 25294
rect 35812 25228 35924 25284
rect 35756 25218 35812 25228
rect 35868 24948 35924 25228
rect 35980 25282 36484 25284
rect 35980 25230 35982 25282
rect 36034 25230 36484 25282
rect 35980 25228 36484 25230
rect 35980 25218 36036 25228
rect 36428 25060 36484 25228
rect 39788 25282 39844 25294
rect 39788 25230 39790 25282
rect 39842 25230 39844 25282
rect 36428 25004 36708 25060
rect 35980 24948 36036 24958
rect 35868 24946 36036 24948
rect 35868 24894 35982 24946
rect 36034 24894 36036 24946
rect 35868 24892 36036 24894
rect 35980 24882 36036 24892
rect 36652 24946 36708 25004
rect 36652 24894 36654 24946
rect 36706 24894 36708 24946
rect 36652 24882 36708 24894
rect 39788 24948 39844 25230
rect 39788 24882 39844 24892
rect 36204 24836 36260 24846
rect 36204 24742 36260 24780
rect 35644 24670 35646 24722
rect 35698 24670 35700 24722
rect 35420 24610 35476 24622
rect 35420 24558 35422 24610
rect 35474 24558 35476 24610
rect 35420 24500 35476 24558
rect 35644 24612 35700 24670
rect 36316 24724 36372 24734
rect 36316 24630 36372 24668
rect 35644 24546 35700 24556
rect 36764 24612 36820 24622
rect 37212 24612 37268 24622
rect 36764 24610 37268 24612
rect 36764 24558 36766 24610
rect 36818 24558 37214 24610
rect 37266 24558 37268 24610
rect 36764 24556 37268 24558
rect 35420 24434 35476 24444
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35420 23940 35476 23950
rect 34636 23938 34916 23940
rect 34636 23886 34638 23938
rect 34690 23886 34916 23938
rect 34636 23884 34916 23886
rect 34636 23874 34692 23884
rect 33516 22306 33572 22316
rect 33852 23548 34132 23604
rect 33404 22260 33460 22270
rect 33404 22166 33460 22204
rect 33852 22260 33908 23548
rect 34860 23378 34916 23884
rect 35420 23846 35476 23884
rect 35868 23940 35924 23950
rect 35868 23846 35924 23884
rect 36764 23604 36820 24556
rect 37212 24546 37268 24556
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 39004 23940 39060 23950
rect 39004 23846 39060 23884
rect 36764 23538 36820 23548
rect 38332 23604 38388 23614
rect 34860 23326 34862 23378
rect 34914 23326 34916 23378
rect 34860 23314 34916 23326
rect 34076 23268 34132 23278
rect 34076 23174 34132 23212
rect 34636 23268 34692 23278
rect 33852 22166 33908 22204
rect 33964 23154 34020 23166
rect 33964 23102 33966 23154
rect 34018 23102 34020 23154
rect 33964 23044 34020 23102
rect 34524 23154 34580 23166
rect 34524 23102 34526 23154
rect 34578 23102 34580 23154
rect 34524 23044 34580 23102
rect 33964 22988 34580 23044
rect 33964 22260 34020 22988
rect 34636 22932 34692 23212
rect 34412 22876 34692 22932
rect 34412 22594 34468 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34412 22542 34414 22594
rect 34466 22542 34468 22594
rect 34412 22530 34468 22542
rect 35084 22484 35140 22494
rect 34972 22372 35028 22382
rect 34972 22278 35028 22316
rect 33964 22258 34132 22260
rect 33964 22206 33966 22258
rect 34018 22206 34132 22258
rect 33964 22204 34132 22206
rect 33964 22194 34020 22204
rect 33180 21970 33236 21980
rect 33292 22146 33348 22158
rect 33292 22094 33294 22146
rect 33346 22094 33348 22146
rect 33292 21924 33348 22094
rect 33628 22146 33684 22158
rect 33628 22094 33630 22146
rect 33682 22094 33684 22146
rect 33628 22036 33684 22094
rect 33292 21858 33348 21868
rect 33404 21980 33684 22036
rect 32732 21746 32788 21756
rect 32508 21588 32564 21626
rect 32508 21522 32564 21532
rect 32508 21364 32564 21374
rect 33068 21364 33124 21374
rect 32508 21362 33124 21364
rect 32508 21310 32510 21362
rect 32562 21310 33070 21362
rect 33122 21310 33124 21362
rect 32508 21308 33124 21310
rect 32508 21298 32564 21308
rect 33068 21298 33124 21308
rect 33292 21364 33348 21374
rect 33292 21270 33348 21308
rect 33404 21140 33460 21980
rect 33740 21812 33796 21822
rect 33740 21718 33796 21756
rect 33628 21700 33684 21710
rect 33628 21588 33684 21644
rect 33852 21700 33908 21710
rect 33852 21606 33908 21644
rect 33964 21588 34020 21598
rect 33628 21586 33796 21588
rect 33628 21534 33630 21586
rect 33682 21534 33796 21586
rect 33628 21532 33796 21534
rect 33628 21522 33684 21532
rect 33068 21084 33460 21140
rect 33068 21026 33124 21084
rect 33068 20974 33070 21026
rect 33122 20974 33124 21026
rect 33068 20962 33124 20974
rect 33628 20916 33684 20926
rect 33628 20822 33684 20860
rect 32844 20804 32900 20814
rect 32844 20710 32900 20748
rect 33740 20802 33796 21532
rect 33964 21494 34020 21532
rect 33964 21028 34020 21038
rect 34076 21028 34132 22204
rect 34524 22258 34580 22270
rect 34524 22206 34526 22258
rect 34578 22206 34580 22258
rect 34412 22148 34468 22158
rect 33964 21026 34132 21028
rect 33964 20974 33966 21026
rect 34018 20974 34132 21026
rect 33964 20972 34132 20974
rect 34188 22146 34468 22148
rect 34188 22094 34414 22146
rect 34466 22094 34468 22146
rect 34188 22092 34468 22094
rect 33964 20962 34020 20972
rect 34188 20916 34244 22092
rect 34412 22082 34468 22092
rect 34524 21812 34580 22206
rect 33740 20750 33742 20802
rect 33794 20750 33796 20802
rect 33740 20692 33796 20750
rect 32284 19954 32340 19964
rect 32396 20578 32452 20590
rect 32396 20526 32398 20578
rect 32450 20526 32452 20578
rect 32396 19460 32452 20526
rect 32508 20578 32564 20590
rect 32508 20526 32510 20578
rect 32562 20526 32564 20578
rect 32508 20356 32564 20526
rect 32620 20580 32676 20590
rect 32620 20486 32676 20524
rect 32508 20300 33460 20356
rect 33404 20130 33460 20300
rect 33740 20244 33796 20636
rect 34076 20860 34244 20916
rect 34300 21756 34580 21812
rect 34076 20244 34132 20860
rect 34300 20804 34356 21756
rect 34636 21700 34692 21710
rect 34692 21644 34916 21700
rect 34636 21634 34692 21644
rect 34524 21586 34580 21598
rect 34524 21534 34526 21586
rect 34578 21534 34580 21586
rect 33404 20078 33406 20130
rect 33458 20078 33460 20130
rect 33404 20066 33460 20078
rect 33516 20188 33796 20244
rect 33852 20188 34132 20244
rect 34188 20748 34356 20804
rect 34412 20916 34468 20926
rect 34412 20802 34468 20860
rect 34412 20750 34414 20802
rect 34466 20750 34468 20802
rect 32508 19906 32564 19918
rect 32508 19854 32510 19906
rect 32562 19854 32564 19906
rect 32508 19796 32564 19854
rect 32508 19730 32564 19740
rect 32396 19404 33236 19460
rect 32620 19124 32676 19134
rect 32620 19030 32676 19068
rect 32060 18958 32062 19010
rect 32114 18958 32116 19010
rect 32060 17108 32116 18958
rect 32732 19010 32788 19022
rect 32732 18958 32734 19010
rect 32786 18958 32788 19010
rect 32732 18900 32788 18958
rect 32172 18340 32228 18350
rect 32172 18246 32228 18284
rect 32620 18228 32676 18238
rect 32732 18228 32788 18844
rect 33180 18450 33236 19404
rect 33516 18900 33572 20188
rect 33628 20018 33684 20030
rect 33628 19966 33630 20018
rect 33682 19966 33684 20018
rect 33628 19572 33684 19966
rect 33628 19506 33684 19516
rect 33516 18834 33572 18844
rect 33740 19234 33796 19246
rect 33740 19182 33742 19234
rect 33794 19182 33796 19234
rect 33180 18398 33182 18450
rect 33234 18398 33236 18450
rect 33180 18386 33236 18398
rect 33740 18340 33796 19182
rect 33740 18274 33796 18284
rect 33852 18450 33908 20188
rect 34188 20132 34244 20748
rect 34412 20244 34468 20750
rect 34524 20580 34580 21534
rect 34860 21586 34916 21644
rect 34860 21534 34862 21586
rect 34914 21534 34916 21586
rect 34860 21522 34916 21534
rect 35084 21364 35140 22428
rect 35868 22484 35924 22494
rect 35868 22390 35924 22428
rect 35420 22260 35476 22270
rect 35420 22166 35476 22204
rect 37436 21812 37492 21822
rect 38220 21812 38276 21822
rect 37436 21810 38276 21812
rect 37436 21758 37438 21810
rect 37490 21758 38222 21810
rect 38274 21758 38276 21810
rect 37436 21756 38276 21758
rect 37436 21746 37492 21756
rect 38220 21746 38276 21756
rect 38332 21698 38388 23548
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 39004 23436 39396 23492
rect 39004 23378 39060 23436
rect 39004 23326 39006 23378
rect 39058 23326 39060 23378
rect 39004 23314 39060 23326
rect 39228 23266 39284 23278
rect 39228 23214 39230 23266
rect 39282 23214 39284 23266
rect 38556 23044 38612 23054
rect 38556 22950 38612 22988
rect 38332 21646 38334 21698
rect 38386 21646 38388 21698
rect 35084 21298 35140 21308
rect 37996 21588 38052 21598
rect 38332 21588 38388 21646
rect 39116 22370 39172 22382
rect 39116 22318 39118 22370
rect 39170 22318 39172 22370
rect 37996 21362 38052 21532
rect 37996 21310 37998 21362
rect 38050 21310 38052 21362
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35420 21028 35476 21038
rect 35420 20934 35476 20972
rect 37996 21028 38052 21310
rect 37996 20962 38052 20972
rect 38108 21532 38388 21588
rect 39004 21586 39060 21598
rect 39004 21534 39006 21586
rect 39058 21534 39060 21586
rect 35532 20916 35588 20926
rect 35532 20822 35588 20860
rect 35084 20804 35140 20814
rect 35084 20710 35140 20748
rect 35196 20802 35252 20814
rect 37884 20804 37940 20814
rect 38108 20804 38164 21532
rect 35196 20750 35198 20802
rect 35250 20750 35252 20802
rect 35196 20692 35252 20750
rect 35196 20626 35252 20636
rect 37548 20802 38164 20804
rect 37548 20750 37886 20802
rect 37938 20750 38164 20802
rect 37548 20748 38164 20750
rect 34524 20514 34580 20524
rect 34972 20580 35028 20590
rect 34076 20020 34132 20030
rect 34188 20020 34244 20076
rect 34076 20018 34244 20020
rect 34076 19966 34078 20018
rect 34130 19966 34244 20018
rect 34076 19964 34244 19966
rect 34076 19954 34132 19964
rect 34188 19346 34244 19964
rect 34300 20188 34468 20244
rect 34300 19458 34356 20188
rect 34972 20018 35028 20524
rect 36092 20580 36148 20590
rect 36092 20486 36148 20524
rect 35308 20020 35364 20030
rect 34972 19966 34974 20018
rect 35026 19966 35028 20018
rect 34412 19796 34468 19806
rect 34412 19794 34804 19796
rect 34412 19742 34414 19794
rect 34466 19742 34804 19794
rect 34412 19740 34804 19742
rect 34412 19730 34468 19740
rect 34300 19406 34302 19458
rect 34354 19406 34356 19458
rect 34300 19394 34356 19406
rect 34188 19294 34190 19346
rect 34242 19294 34244 19346
rect 34188 19282 34244 19294
rect 34748 19234 34804 19740
rect 34748 19182 34750 19234
rect 34802 19182 34804 19234
rect 34748 19170 34804 19182
rect 33852 18398 33854 18450
rect 33906 18398 33908 18450
rect 32620 18226 32788 18228
rect 32620 18174 32622 18226
rect 32674 18174 32788 18226
rect 32620 18172 32788 18174
rect 33852 18228 33908 18398
rect 32620 18162 32676 18172
rect 33852 17666 33908 18172
rect 34076 19124 34132 19134
rect 34076 18338 34132 19068
rect 34076 18286 34078 18338
rect 34130 18286 34132 18338
rect 34076 17892 34132 18286
rect 34636 18340 34692 18350
rect 34748 18340 34804 18350
rect 34636 18338 34748 18340
rect 34636 18286 34638 18338
rect 34690 18286 34748 18338
rect 34636 18284 34748 18286
rect 34636 18274 34692 18284
rect 34524 18228 34580 18238
rect 34524 18134 34580 18172
rect 34076 17836 34468 17892
rect 33852 17614 33854 17666
rect 33906 17614 33908 17666
rect 33852 17602 33908 17614
rect 34300 17666 34356 17678
rect 34300 17614 34302 17666
rect 34354 17614 34356 17666
rect 32844 17444 32900 17454
rect 33404 17444 33460 17454
rect 32844 17350 32900 17388
rect 33180 17442 33460 17444
rect 33180 17390 33406 17442
rect 33458 17390 33460 17442
rect 33180 17388 33460 17390
rect 33180 17108 33236 17388
rect 33404 17378 33460 17388
rect 33628 17442 33684 17454
rect 33628 17390 33630 17442
rect 33682 17390 33684 17442
rect 33628 17108 33684 17390
rect 32060 17042 32116 17052
rect 32620 17106 33236 17108
rect 32620 17054 33182 17106
rect 33234 17054 33236 17106
rect 32620 17052 33236 17054
rect 32060 16212 32116 16222
rect 31948 16210 32116 16212
rect 31948 16158 32062 16210
rect 32114 16158 32116 16210
rect 31948 16156 32116 16158
rect 31948 15426 32004 16156
rect 32060 16146 32116 16156
rect 32172 16044 32564 16100
rect 31948 15374 31950 15426
rect 32002 15374 32004 15426
rect 31948 15362 32004 15374
rect 32060 15874 32116 15886
rect 32060 15822 32062 15874
rect 32114 15822 32116 15874
rect 32060 15764 32116 15822
rect 32172 15874 32228 16044
rect 32172 15822 32174 15874
rect 32226 15822 32228 15874
rect 32172 15810 32228 15822
rect 32396 15876 32452 15886
rect 32396 15782 32452 15820
rect 32508 15764 32564 16044
rect 32620 16098 32676 17052
rect 33180 17042 33236 17052
rect 33516 17052 33684 17108
rect 33740 17442 33796 17454
rect 33740 17390 33742 17442
rect 33794 17390 33796 17442
rect 33740 17108 33796 17390
rect 33740 17052 34132 17108
rect 33292 16996 33348 17006
rect 33180 16660 33236 16670
rect 33180 16566 33236 16604
rect 33292 16212 33348 16940
rect 33292 16146 33348 16156
rect 32620 16046 32622 16098
rect 32674 16046 32676 16098
rect 32620 16034 32676 16046
rect 32956 16098 33012 16110
rect 32956 16046 32958 16098
rect 33010 16046 33012 16098
rect 32956 15764 33012 16046
rect 33292 15988 33348 15998
rect 33292 15894 33348 15932
rect 32508 15708 32788 15764
rect 32060 15316 32116 15708
rect 32284 15652 32340 15662
rect 32060 15250 32116 15260
rect 32172 15540 32228 15550
rect 32172 15148 32228 15484
rect 31500 15138 31556 15148
rect 31612 15092 31892 15148
rect 32060 15092 32228 15148
rect 31500 14868 31556 14878
rect 31500 13300 31556 14812
rect 31612 13748 31668 15092
rect 32060 15090 32116 15092
rect 32060 15038 32062 15090
rect 32114 15038 32116 15090
rect 32060 15026 32116 15038
rect 32284 14756 32340 15596
rect 32620 15316 32676 15326
rect 32508 15260 32620 15316
rect 32508 15202 32564 15260
rect 32620 15250 32676 15260
rect 32508 15150 32510 15202
rect 32562 15150 32564 15202
rect 32508 15138 32564 15150
rect 32732 15148 32788 15708
rect 32956 15698 33012 15708
rect 33180 15874 33236 15886
rect 33180 15822 33182 15874
rect 33234 15822 33236 15874
rect 33180 15540 33236 15822
rect 33404 15876 33460 15886
rect 33516 15876 33572 17052
rect 33628 16884 33684 16894
rect 33628 16790 33684 16828
rect 34076 16882 34132 17052
rect 34076 16830 34078 16882
rect 34130 16830 34132 16882
rect 34076 16818 34132 16830
rect 34188 16996 34244 17006
rect 33628 16156 34132 16212
rect 33628 16098 33684 16156
rect 33628 16046 33630 16098
rect 33682 16046 33684 16098
rect 33628 16034 33684 16046
rect 33964 15988 34020 15998
rect 33740 15986 34020 15988
rect 33740 15934 33966 15986
rect 34018 15934 34020 15986
rect 33740 15932 34020 15934
rect 33740 15876 33796 15932
rect 33516 15820 33796 15876
rect 33404 15782 33460 15820
rect 31948 14700 32340 14756
rect 32620 15092 32788 15148
rect 32844 15484 33236 15540
rect 32620 14980 32676 15092
rect 31948 14642 32004 14700
rect 31948 14590 31950 14642
rect 32002 14590 32004 14642
rect 31948 14578 32004 14590
rect 32508 13860 32564 13870
rect 32620 13860 32676 14924
rect 32564 13804 32676 13860
rect 32732 14418 32788 14430
rect 32732 14366 32734 14418
rect 32786 14366 32788 14418
rect 32508 13766 32564 13804
rect 31612 13654 31668 13692
rect 32060 13746 32116 13758
rect 32284 13748 32340 13758
rect 32060 13694 32062 13746
rect 32114 13694 32116 13746
rect 32060 13636 32116 13694
rect 31948 13580 32060 13636
rect 31948 13524 32004 13580
rect 32060 13570 32116 13580
rect 32172 13692 32284 13748
rect 31836 13468 32004 13524
rect 31500 13244 31668 13300
rect 31500 13076 31556 13086
rect 31388 13074 31556 13076
rect 31388 13022 31502 13074
rect 31554 13022 31556 13074
rect 31388 13020 31556 13022
rect 31164 11396 31220 11406
rect 31164 11302 31220 11340
rect 31052 11190 31108 11228
rect 31276 11284 31332 11322
rect 31276 11218 31332 11228
rect 30940 10770 30996 10780
rect 31276 10836 31332 10846
rect 31276 10742 31332 10780
rect 30716 9650 30772 9660
rect 30940 10498 30996 10510
rect 30940 10446 30942 10498
rect 30994 10446 30996 10498
rect 30492 9602 30548 9614
rect 30492 9550 30494 9602
rect 30546 9550 30548 9602
rect 30380 9268 30436 9278
rect 30380 9174 30436 9212
rect 30268 9154 30324 9166
rect 30268 9102 30270 9154
rect 30322 9102 30324 9154
rect 30268 8820 30324 9102
rect 30492 9156 30548 9550
rect 30828 9604 30884 9614
rect 30828 9510 30884 9548
rect 30940 9492 30996 10446
rect 31388 9828 31444 13020
rect 31500 13010 31556 13020
rect 31612 11788 31668 13244
rect 31836 13186 31892 13468
rect 32172 13412 32228 13692
rect 31836 13134 31838 13186
rect 31890 13134 31892 13186
rect 31836 13122 31892 13134
rect 31948 13356 32228 13412
rect 31948 13074 32004 13356
rect 31948 13022 31950 13074
rect 32002 13022 32004 13074
rect 31948 13010 32004 13022
rect 32284 12404 32340 13692
rect 32732 13748 32788 14366
rect 32732 13682 32788 13692
rect 32844 14418 32900 15484
rect 33740 15428 33796 15820
rect 33964 15876 34020 15932
rect 34076 15988 34132 16156
rect 34188 15988 34244 16940
rect 34300 16098 34356 17614
rect 34300 16046 34302 16098
rect 34354 16046 34356 16098
rect 34300 16034 34356 16046
rect 34076 15986 34244 15988
rect 34076 15934 34078 15986
rect 34130 15934 34244 15986
rect 34076 15932 34244 15934
rect 34076 15922 34132 15932
rect 33964 15810 34020 15820
rect 34412 15764 34468 17836
rect 34636 17780 34692 17790
rect 34636 17686 34692 17724
rect 34524 17444 34580 17454
rect 34524 17350 34580 17388
rect 34636 16324 34692 16334
rect 34636 16230 34692 16268
rect 34524 15988 34580 15998
rect 34524 15894 34580 15932
rect 34748 15764 34804 18284
rect 34972 18340 35028 19966
rect 35084 20018 35364 20020
rect 35084 19966 35310 20018
rect 35362 19966 35364 20018
rect 35084 19964 35364 19966
rect 35084 19122 35140 19964
rect 35308 19954 35364 19964
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35532 19460 35588 19470
rect 35532 19346 35588 19404
rect 35532 19294 35534 19346
rect 35586 19294 35588 19346
rect 35532 19282 35588 19294
rect 37212 19348 37268 19358
rect 37548 19348 37604 20748
rect 37884 20738 37940 20748
rect 39004 20468 39060 21534
rect 39116 21588 39172 22318
rect 39116 21522 39172 21532
rect 39004 20402 39060 20412
rect 37660 20130 37716 20142
rect 37660 20078 37662 20130
rect 37714 20078 37716 20130
rect 37660 19458 37716 20078
rect 38444 20132 38500 20142
rect 38444 20020 38500 20076
rect 39228 20132 39284 23214
rect 39340 23156 39396 23436
rect 39900 23266 39956 23278
rect 39900 23214 39902 23266
rect 39954 23214 39956 23266
rect 39564 23156 39620 23166
rect 39340 23154 39620 23156
rect 39340 23102 39566 23154
rect 39618 23102 39620 23154
rect 39340 23100 39620 23102
rect 39564 21588 39620 23100
rect 39900 22148 39956 23214
rect 40236 23154 40292 23166
rect 40236 23102 40238 23154
rect 40290 23102 40292 23154
rect 40236 22932 40292 23102
rect 40236 22866 40292 22876
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 39900 22082 39956 22092
rect 39564 21522 39620 21532
rect 40124 21474 40180 21486
rect 40124 21422 40126 21474
rect 40178 21422 40180 21474
rect 40124 20916 40180 21422
rect 40124 20850 40180 20860
rect 40236 20690 40292 20702
rect 40236 20638 40238 20690
rect 40290 20638 40292 20690
rect 39676 20578 39732 20590
rect 39676 20526 39678 20578
rect 39730 20526 39732 20578
rect 39676 20244 39732 20526
rect 39676 20178 39732 20188
rect 39900 20578 39956 20590
rect 39900 20526 39902 20578
rect 39954 20526 39956 20578
rect 39228 20066 39284 20076
rect 39004 20020 39060 20030
rect 38444 20018 39060 20020
rect 38444 19966 39006 20018
rect 39058 19966 39060 20018
rect 38444 19964 39060 19966
rect 39004 19954 39060 19964
rect 37660 19406 37662 19458
rect 37714 19406 37716 19458
rect 37660 19394 37716 19406
rect 37212 19346 37604 19348
rect 37212 19294 37214 19346
rect 37266 19294 37550 19346
rect 37602 19294 37604 19346
rect 37212 19292 37604 19294
rect 37212 19282 37268 19292
rect 35084 19070 35086 19122
rect 35138 19070 35140 19122
rect 35084 19058 35140 19070
rect 35980 19010 36036 19022
rect 35980 18958 35982 19010
rect 36034 18958 36036 19010
rect 35084 18340 35140 18350
rect 34972 18338 35140 18340
rect 34972 18286 35086 18338
rect 35138 18286 35140 18338
rect 34972 18284 35140 18286
rect 34972 17556 35028 18284
rect 35084 18274 35140 18284
rect 35532 18340 35588 18350
rect 35980 18340 36036 18958
rect 35588 18284 36036 18340
rect 35532 18246 35588 18284
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35980 17780 36036 17790
rect 36036 17724 36148 17780
rect 35980 17686 36036 17724
rect 34860 16884 34916 16894
rect 34972 16884 35028 17500
rect 35532 17556 35588 17566
rect 35532 17462 35588 17500
rect 34916 16828 35028 16884
rect 34860 16818 34916 16828
rect 34412 15698 34468 15708
rect 34524 15708 34804 15764
rect 34860 15764 34916 15774
rect 33740 15362 33796 15372
rect 33292 15314 33348 15326
rect 33292 15262 33294 15314
rect 33346 15262 33348 15314
rect 33180 15092 33236 15102
rect 32844 14366 32846 14418
rect 32898 14366 32900 14418
rect 32396 13634 32452 13646
rect 32396 13582 32398 13634
rect 32450 13582 32452 13634
rect 32396 13188 32452 13582
rect 32844 13636 32900 14366
rect 32956 14420 33012 14430
rect 32956 14326 33012 14364
rect 33068 13972 33124 13982
rect 33068 13858 33124 13916
rect 33180 13970 33236 15036
rect 33292 14980 33348 15262
rect 33628 15316 33684 15326
rect 33628 15222 33684 15260
rect 33852 15316 33908 15326
rect 34076 15316 34132 15326
rect 33852 15314 34132 15316
rect 33852 15262 33854 15314
rect 33906 15262 34078 15314
rect 34130 15262 34132 15314
rect 33852 15260 34132 15262
rect 33292 14914 33348 14924
rect 33404 15202 33460 15214
rect 33404 15150 33406 15202
rect 33458 15150 33460 15202
rect 33404 14532 33460 15150
rect 33852 15148 33908 15260
rect 34076 15250 34132 15260
rect 34412 15314 34468 15326
rect 34412 15262 34414 15314
rect 34466 15262 34468 15314
rect 34412 15148 34468 15262
rect 33180 13918 33182 13970
rect 33234 13918 33236 13970
rect 33180 13906 33236 13918
rect 33292 14476 33460 14532
rect 33628 15092 33908 15148
rect 34188 15092 34468 15148
rect 33068 13806 33070 13858
rect 33122 13806 33124 13858
rect 33068 13794 33124 13806
rect 32844 13570 32900 13580
rect 32508 13188 32564 13198
rect 32396 13186 32564 13188
rect 32396 13134 32510 13186
rect 32562 13134 32564 13186
rect 32396 13132 32564 13134
rect 32508 13122 32564 13132
rect 32732 13188 32788 13198
rect 32732 13094 32788 13132
rect 33068 12962 33124 12974
rect 33068 12910 33070 12962
rect 33122 12910 33124 12962
rect 33068 12852 33124 12910
rect 33180 12964 33236 12974
rect 33292 12964 33348 14476
rect 33404 14308 33460 14318
rect 33404 14306 33572 14308
rect 33404 14254 33406 14306
rect 33458 14254 33572 14306
rect 33404 14252 33572 14254
rect 33404 14242 33460 14252
rect 33180 12962 33348 12964
rect 33180 12910 33182 12962
rect 33234 12910 33348 12962
rect 33180 12908 33348 12910
rect 33404 13746 33460 13758
rect 33404 13694 33406 13746
rect 33458 13694 33460 13746
rect 33404 12962 33460 13694
rect 33516 13188 33572 14252
rect 33628 13858 33684 15092
rect 34188 14530 34244 15092
rect 34188 14478 34190 14530
rect 34242 14478 34244 14530
rect 34188 14420 34244 14478
rect 34188 13972 34244 14364
rect 34188 13906 34244 13916
rect 34524 13860 34580 15708
rect 34636 15540 34692 15550
rect 34860 15540 34916 15708
rect 34636 15538 34916 15540
rect 34636 15486 34638 15538
rect 34690 15486 34916 15538
rect 34636 15484 34916 15486
rect 34636 15316 34692 15484
rect 34636 15250 34692 15260
rect 34972 15148 35028 16828
rect 35084 17442 35140 17454
rect 35084 17390 35086 17442
rect 35138 17390 35140 17442
rect 35084 15876 35140 17390
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35532 16212 35588 16222
rect 35532 16118 35588 16156
rect 36092 16210 36148 17724
rect 36428 16996 36484 17006
rect 36204 16994 36484 16996
rect 36204 16942 36430 16994
rect 36482 16942 36484 16994
rect 36204 16940 36484 16942
rect 36204 16322 36260 16940
rect 36428 16930 36484 16940
rect 37212 16996 37268 17006
rect 37212 16902 37268 16940
rect 36204 16270 36206 16322
rect 36258 16270 36260 16322
rect 36204 16258 36260 16270
rect 36092 16158 36094 16210
rect 36146 16158 36148 16210
rect 35084 15782 35140 15820
rect 35532 15876 35588 15886
rect 35532 15538 35588 15820
rect 35532 15486 35534 15538
rect 35586 15486 35588 15538
rect 35532 15474 35588 15486
rect 36092 15538 36148 16158
rect 36092 15486 36094 15538
rect 36146 15486 36148 15538
rect 36092 15474 36148 15486
rect 35084 15202 35140 15214
rect 35084 15150 35086 15202
rect 35138 15150 35140 15202
rect 35084 15148 35140 15150
rect 34748 15092 34804 15102
rect 34748 14998 34804 15036
rect 34860 15092 35140 15148
rect 35756 15092 35812 15102
rect 33628 13806 33630 13858
rect 33682 13806 33684 13858
rect 33628 13794 33684 13806
rect 34412 13804 34580 13860
rect 34636 14980 34692 14990
rect 34636 14642 34692 14924
rect 34636 14590 34638 14642
rect 34690 14590 34692 14642
rect 34076 13748 34132 13758
rect 34412 13748 34468 13804
rect 33964 13746 34468 13748
rect 33964 13694 34078 13746
rect 34130 13694 34468 13746
rect 33964 13692 34468 13694
rect 33572 13132 33684 13188
rect 33516 13122 33572 13132
rect 33404 12910 33406 12962
rect 33458 12910 33460 12962
rect 33180 12898 33236 12908
rect 33404 12898 33460 12910
rect 32396 12404 32452 12414
rect 32284 12402 32452 12404
rect 32284 12350 32398 12402
rect 32450 12350 32452 12402
rect 32284 12348 32452 12350
rect 32396 12338 32452 12348
rect 33068 12178 33124 12796
rect 33068 12126 33070 12178
rect 33122 12126 33124 12178
rect 33068 12114 33124 12126
rect 33292 12738 33348 12750
rect 33292 12686 33294 12738
rect 33346 12686 33348 12738
rect 30492 9100 30884 9156
rect 30268 8754 30324 8764
rect 30156 8318 30158 8370
rect 30210 8318 30212 8370
rect 30156 8306 30212 8318
rect 30604 8372 30660 8382
rect 30604 8278 30660 8316
rect 29708 8206 29710 8258
rect 29762 8206 29764 8258
rect 29708 8194 29764 8206
rect 28476 8094 28478 8146
rect 28530 8094 28532 8146
rect 28476 8082 28532 8094
rect 28588 8146 28644 8158
rect 28588 8094 28590 8146
rect 28642 8094 28644 8146
rect 28588 8036 28644 8094
rect 29260 8036 29316 8046
rect 28588 8034 29316 8036
rect 28588 7982 29262 8034
rect 29314 7982 29316 8034
rect 28588 7980 29316 7982
rect 29260 7970 29316 7980
rect 27916 7698 28196 7700
rect 27916 7646 27918 7698
rect 27970 7646 28196 7698
rect 27916 7644 28196 7646
rect 27916 7634 27972 7644
rect 28700 7588 28756 7598
rect 28700 7494 28756 7532
rect 30828 7476 30884 9100
rect 30940 8930 30996 9436
rect 30940 8878 30942 8930
rect 30994 8878 30996 8930
rect 30940 8372 30996 8878
rect 31276 9772 31444 9828
rect 31500 11732 31668 11788
rect 32060 11956 32116 11966
rect 33292 11956 33348 12686
rect 33628 12404 33684 13132
rect 33628 12178 33684 12348
rect 33740 12292 33796 12302
rect 33740 12198 33796 12236
rect 33628 12126 33630 12178
rect 33682 12126 33684 12178
rect 33628 12114 33684 12126
rect 31500 10834 31556 11732
rect 31836 11396 31892 11406
rect 31500 10782 31502 10834
rect 31554 10782 31556 10834
rect 30940 8306 30996 8316
rect 31164 8372 31220 8382
rect 31164 8278 31220 8316
rect 31276 8260 31332 9772
rect 31500 9716 31556 10782
rect 31724 11282 31780 11294
rect 31724 11230 31726 11282
rect 31778 11230 31780 11282
rect 31612 10724 31668 10734
rect 31724 10724 31780 11230
rect 31668 10668 31780 10724
rect 31612 10630 31668 10668
rect 31500 9650 31556 9660
rect 31388 9602 31444 9614
rect 31388 9550 31390 9602
rect 31442 9550 31444 9602
rect 31388 9492 31444 9550
rect 31388 9426 31444 9436
rect 31500 9156 31556 9166
rect 31500 9062 31556 9100
rect 31612 9044 31668 9054
rect 31612 8950 31668 8988
rect 31836 8932 31892 11340
rect 32060 11394 32116 11900
rect 32060 11342 32062 11394
rect 32114 11342 32116 11394
rect 32060 11330 32116 11342
rect 32732 11900 33348 11956
rect 33964 11956 34020 13692
rect 34076 13682 34132 13692
rect 34524 13636 34580 13646
rect 34076 13524 34132 13534
rect 34076 12962 34132 13468
rect 34188 13188 34244 13198
rect 34188 13074 34244 13132
rect 34188 13022 34190 13074
rect 34242 13022 34244 13074
rect 34188 13010 34244 13022
rect 34076 12910 34078 12962
rect 34130 12910 34132 12962
rect 34076 12898 34132 12910
rect 34524 12852 34580 13580
rect 34524 12786 34580 12796
rect 34188 12740 34244 12750
rect 32732 11282 32788 11900
rect 33964 11890 34020 11900
rect 34076 12292 34132 12302
rect 34076 12066 34132 12236
rect 34076 12014 34078 12066
rect 34130 12014 34132 12066
rect 34076 11844 34132 12014
rect 34076 11778 34132 11788
rect 33404 11508 33460 11518
rect 32844 11396 32900 11406
rect 32844 11394 33124 11396
rect 32844 11342 32846 11394
rect 32898 11342 33124 11394
rect 32844 11340 33124 11342
rect 32844 11330 32900 11340
rect 32732 11230 32734 11282
rect 32786 11230 32788 11282
rect 32732 11218 32788 11230
rect 32060 10722 32116 10734
rect 32060 10670 32062 10722
rect 32114 10670 32116 10722
rect 32060 10052 32116 10670
rect 33068 10722 33124 11340
rect 33404 11394 33460 11452
rect 33404 11342 33406 11394
rect 33458 11342 33460 11394
rect 33404 11330 33460 11342
rect 33740 11396 33796 11406
rect 34188 11396 34244 12684
rect 34300 12740 34356 12750
rect 34636 12740 34692 14590
rect 34860 14308 34916 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 34860 13746 34916 14252
rect 35644 14306 35700 14318
rect 35644 14254 35646 14306
rect 35698 14254 35700 14306
rect 34860 13694 34862 13746
rect 34914 13694 34916 13746
rect 34748 12964 34804 12974
rect 34748 12870 34804 12908
rect 34300 12738 34468 12740
rect 34300 12686 34302 12738
rect 34354 12686 34468 12738
rect 34300 12684 34468 12686
rect 34300 12674 34356 12684
rect 33068 10670 33070 10722
rect 33122 10670 33124 10722
rect 33068 10658 33124 10670
rect 32284 10610 32340 10622
rect 32284 10558 32286 10610
rect 32338 10558 32340 10610
rect 32284 10388 32340 10558
rect 32508 10612 32564 10622
rect 32508 10610 33012 10612
rect 32508 10558 32510 10610
rect 32562 10558 33012 10610
rect 32508 10556 33012 10558
rect 32508 10546 32564 10556
rect 32284 10322 32340 10332
rect 32396 10498 32452 10510
rect 32396 10446 32398 10498
rect 32450 10446 32452 10498
rect 32060 9986 32116 9996
rect 32284 9716 32340 9726
rect 31948 9604 32004 9614
rect 31948 9266 32004 9548
rect 31948 9214 31950 9266
rect 32002 9214 32004 9266
rect 31948 9202 32004 9214
rect 32172 9268 32228 9278
rect 32284 9268 32340 9660
rect 32396 9380 32452 10446
rect 32844 9826 32900 9838
rect 32844 9774 32846 9826
rect 32898 9774 32900 9826
rect 32844 9716 32900 9774
rect 32956 9716 33012 10556
rect 33740 10610 33796 11340
rect 34076 11394 34244 11396
rect 34076 11342 34190 11394
rect 34242 11342 34244 11394
rect 34076 11340 34244 11342
rect 33964 11284 34020 11294
rect 33964 11170 34020 11228
rect 33964 11118 33966 11170
rect 34018 11118 34020 11170
rect 33964 11106 34020 11118
rect 33740 10558 33742 10610
rect 33794 10558 33796 10610
rect 33740 10546 33796 10558
rect 33964 10612 34020 10622
rect 34076 10612 34132 11340
rect 34188 11330 34244 11340
rect 34300 11172 34356 11182
rect 34300 11078 34356 11116
rect 33964 10610 34132 10612
rect 33964 10558 33966 10610
rect 34018 10558 34132 10610
rect 33964 10556 34132 10558
rect 33964 10546 34020 10556
rect 34300 10388 34356 10398
rect 34412 10388 34468 12684
rect 34636 12674 34692 12684
rect 34524 12404 34580 12414
rect 34524 12310 34580 12348
rect 34748 12180 34804 12190
rect 34636 12068 34692 12078
rect 34636 11974 34692 12012
rect 34524 11396 34580 11406
rect 34524 11302 34580 11340
rect 34748 11394 34804 12124
rect 34748 11342 34750 11394
rect 34802 11342 34804 11394
rect 34356 10332 34468 10388
rect 34300 10322 34356 10332
rect 34636 10052 34692 10062
rect 34636 9958 34692 9996
rect 33516 9940 33572 9950
rect 32956 9660 33460 9716
rect 32844 9650 32900 9660
rect 32396 9324 33236 9380
rect 32172 9266 32284 9268
rect 32172 9214 32174 9266
rect 32226 9214 32284 9266
rect 32172 9212 32284 9214
rect 32060 9044 32116 9054
rect 32060 8950 32116 8988
rect 31836 8866 31892 8876
rect 31500 8820 31556 8830
rect 31500 8726 31556 8764
rect 31724 8372 31780 8382
rect 32172 8372 32228 9212
rect 32284 9174 32340 9212
rect 32620 9044 32676 9054
rect 32620 8950 32676 8988
rect 33068 9042 33124 9054
rect 33068 8990 33070 9042
rect 33122 8990 33124 9042
rect 33068 8932 33124 8990
rect 33068 8866 33124 8876
rect 31780 8370 32228 8372
rect 31780 8318 32174 8370
rect 32226 8318 32228 8370
rect 31780 8316 32228 8318
rect 31724 8278 31780 8316
rect 32172 8306 32228 8316
rect 30940 7476 30996 7486
rect 30828 7474 30996 7476
rect 30828 7422 30942 7474
rect 30994 7422 30996 7474
rect 30828 7420 30996 7422
rect 31276 7476 31332 8204
rect 32620 8260 32676 8270
rect 32620 8166 32676 8204
rect 33068 8260 33124 8270
rect 31948 8148 32004 8158
rect 31836 7588 31892 7598
rect 31836 7494 31892 7532
rect 31948 7588 32004 8092
rect 33068 7700 33124 8204
rect 33180 8258 33236 9324
rect 33404 9266 33460 9660
rect 33404 9214 33406 9266
rect 33458 9214 33460 9266
rect 33404 9202 33460 9214
rect 33404 9044 33460 9054
rect 33516 9044 33572 9884
rect 33964 9828 34020 9838
rect 34748 9828 34804 11342
rect 33964 9714 34020 9772
rect 34636 9772 34804 9828
rect 34860 10610 34916 13694
rect 35532 13746 35588 13758
rect 35532 13694 35534 13746
rect 35586 13694 35588 13746
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35532 13188 35588 13694
rect 35644 13748 35700 14254
rect 35644 13682 35700 13692
rect 35532 13122 35588 13132
rect 35308 12964 35364 12974
rect 35308 12962 35700 12964
rect 35308 12910 35310 12962
rect 35362 12910 35700 12962
rect 35308 12908 35700 12910
rect 35308 12898 35364 12908
rect 34972 12852 35028 12862
rect 34972 12516 35028 12796
rect 35644 12850 35700 12908
rect 35756 12962 35812 15036
rect 36092 14308 36148 14318
rect 36092 14214 36148 14252
rect 37324 13076 37380 19292
rect 37548 19282 37604 19292
rect 39900 19348 39956 20526
rect 40236 20244 40292 20638
rect 40236 20178 40292 20188
rect 40012 19906 40068 19918
rect 40012 19854 40014 19906
rect 40066 19854 40068 19906
rect 40012 19572 40068 19854
rect 40012 19506 40068 19516
rect 39900 19282 39956 19292
rect 40236 19122 40292 19134
rect 40236 19070 40238 19122
rect 40290 19070 40292 19122
rect 39676 19010 39732 19022
rect 39676 18958 39678 19010
rect 39730 18958 39732 19010
rect 39676 18900 39732 18958
rect 39900 19012 39956 19022
rect 39900 18918 39956 18956
rect 39676 18834 39732 18844
rect 40236 18900 40292 19070
rect 40236 18834 40292 18844
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 39116 17666 39172 17678
rect 39116 17614 39118 17666
rect 39170 17614 39172 17666
rect 39004 16882 39060 16894
rect 39004 16830 39006 16882
rect 39058 16830 39060 16882
rect 39004 16324 39060 16830
rect 39004 16258 39060 16268
rect 39004 16100 39060 16110
rect 39004 16006 39060 16044
rect 39116 15540 39172 17614
rect 39788 16882 39844 16894
rect 39788 16830 39790 16882
rect 39842 16830 39844 16882
rect 39788 16212 39844 16830
rect 40012 16884 40068 17726
rect 40012 16818 40068 16828
rect 39788 16146 39844 16156
rect 40124 15986 40180 15998
rect 40124 15934 40126 15986
rect 40178 15934 40180 15986
rect 39116 15474 39172 15484
rect 39228 15764 39284 15774
rect 39004 15314 39060 15326
rect 39004 15262 39006 15314
rect 39058 15262 39060 15314
rect 39004 14756 39060 15262
rect 39004 14690 39060 14700
rect 39228 14642 39284 15708
rect 40124 15540 40180 15934
rect 40124 15474 40180 15484
rect 39788 15202 39844 15214
rect 39788 15150 39790 15202
rect 39842 15150 39844 15202
rect 39788 14868 39844 15150
rect 39788 14802 39844 14812
rect 40348 15202 40404 15214
rect 40348 15150 40350 15202
rect 40402 15150 40404 15202
rect 39228 14590 39230 14642
rect 39282 14590 39284 14642
rect 39228 14578 39284 14590
rect 40236 14532 40292 14542
rect 40348 14532 40404 15150
rect 40236 14530 40404 14532
rect 40236 14478 40238 14530
rect 40290 14478 40404 14530
rect 40236 14476 40404 14478
rect 40236 14196 40292 14476
rect 40236 14130 40292 14140
rect 38556 13972 38612 13982
rect 38556 13878 38612 13916
rect 37772 13858 37828 13870
rect 37772 13806 37774 13858
rect 37826 13806 37828 13858
rect 37772 13186 37828 13806
rect 37772 13134 37774 13186
rect 37826 13134 37828 13186
rect 37772 13122 37828 13134
rect 38668 13748 38724 13758
rect 39004 13748 39060 13758
rect 38724 13746 39060 13748
rect 38724 13694 39006 13746
rect 39058 13694 39060 13746
rect 38724 13692 39060 13694
rect 37660 13076 37716 13086
rect 37324 13074 37716 13076
rect 37324 13022 37326 13074
rect 37378 13022 37662 13074
rect 37714 13022 37716 13074
rect 37324 13020 37716 13022
rect 37324 13010 37380 13020
rect 35756 12910 35758 12962
rect 35810 12910 35812 12962
rect 35756 12898 35812 12910
rect 35980 12964 36036 12974
rect 35980 12870 36036 12908
rect 35644 12798 35646 12850
rect 35698 12798 35700 12850
rect 35644 12786 35700 12798
rect 36316 12850 36372 12862
rect 36316 12798 36318 12850
rect 36370 12798 36372 12850
rect 35084 12740 35140 12750
rect 35420 12740 35476 12750
rect 36204 12740 36260 12750
rect 35084 12738 35252 12740
rect 35084 12686 35086 12738
rect 35138 12686 35252 12738
rect 35084 12684 35252 12686
rect 35084 12674 35140 12684
rect 34972 12460 35140 12516
rect 34972 12292 35028 12302
rect 34972 12198 35028 12236
rect 35084 12068 35140 12460
rect 34972 12012 35140 12068
rect 34972 11396 35028 12012
rect 35196 11956 35252 12684
rect 35420 12738 35588 12740
rect 35420 12686 35422 12738
rect 35474 12686 35588 12738
rect 35420 12684 35588 12686
rect 35420 12674 35476 12684
rect 35532 12292 35588 12684
rect 36204 12646 36260 12684
rect 35980 12404 36036 12414
rect 35532 12236 35700 12292
rect 35196 11890 35252 11900
rect 35532 12066 35588 12078
rect 35532 12014 35534 12066
rect 35586 12014 35588 12066
rect 35532 11956 35588 12014
rect 35532 11890 35588 11900
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35644 11620 35700 12236
rect 34972 11330 35028 11340
rect 35532 11564 35700 11620
rect 35980 12066 36036 12348
rect 35980 12014 35982 12066
rect 36034 12014 36036 12066
rect 35980 11956 36036 12014
rect 35084 11284 35140 11294
rect 35084 11190 35140 11228
rect 35196 11170 35252 11182
rect 35196 11118 35198 11170
rect 35250 11118 35252 11170
rect 35196 10948 35252 11118
rect 35308 11172 35364 11182
rect 35308 11170 35476 11172
rect 35308 11118 35310 11170
rect 35362 11118 35476 11170
rect 35308 11116 35476 11118
rect 35308 11106 35364 11116
rect 35196 10892 35364 10948
rect 34860 10558 34862 10610
rect 34914 10558 34916 10610
rect 33964 9662 33966 9714
rect 34018 9662 34020 9714
rect 33852 9604 33908 9614
rect 33404 9042 33572 9044
rect 33404 8990 33406 9042
rect 33458 8990 33572 9042
rect 33404 8988 33572 8990
rect 33740 9602 33908 9604
rect 33740 9550 33854 9602
rect 33906 9550 33908 9602
rect 33740 9548 33908 9550
rect 33740 9042 33796 9548
rect 33852 9538 33908 9548
rect 33852 9156 33908 9166
rect 33852 9062 33908 9100
rect 33740 8990 33742 9042
rect 33794 8990 33796 9042
rect 33404 8978 33460 8988
rect 33740 8978 33796 8990
rect 33964 9044 34020 9662
rect 34188 9716 34244 9726
rect 34076 9268 34132 9278
rect 34076 9174 34132 9212
rect 34188 9154 34244 9660
rect 34636 9716 34692 9772
rect 34636 9622 34692 9660
rect 34748 9658 34804 9670
rect 34748 9606 34750 9658
rect 34802 9606 34804 9658
rect 34748 9604 34804 9606
rect 34748 9538 34804 9548
rect 34636 9268 34692 9278
rect 34860 9268 34916 10558
rect 35308 10610 35364 10892
rect 35308 10558 35310 10610
rect 35362 10558 35364 10610
rect 35308 10546 35364 10558
rect 35308 10388 35364 10398
rect 35420 10388 35476 11116
rect 35364 10332 35476 10388
rect 35308 10322 35364 10332
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35532 9828 35588 11564
rect 35644 11396 35700 11406
rect 35868 11396 35924 11406
rect 35644 11394 35924 11396
rect 35644 11342 35646 11394
rect 35698 11342 35870 11394
rect 35922 11342 35924 11394
rect 35644 11340 35924 11342
rect 35644 11330 35700 11340
rect 35868 11330 35924 11340
rect 35532 9762 35588 9772
rect 35308 9604 35364 9614
rect 35980 9604 36036 11900
rect 36204 11396 36260 11406
rect 36316 11396 36372 12798
rect 36204 11394 36372 11396
rect 36204 11342 36206 11394
rect 36258 11342 36372 11394
rect 36204 11340 36372 11342
rect 36092 11284 36148 11294
rect 36092 11190 36148 11228
rect 35308 9602 36036 9604
rect 35308 9550 35310 9602
rect 35362 9550 36036 9602
rect 35308 9548 36036 9550
rect 36204 9604 36260 11340
rect 37212 11284 37268 11294
rect 37212 11190 37268 11228
rect 37660 10724 37716 13020
rect 38668 13074 38724 13692
rect 39004 13682 39060 13692
rect 40012 13634 40068 13646
rect 40012 13582 40014 13634
rect 40066 13582 40068 13634
rect 40012 13524 40068 13582
rect 40012 13458 40068 13468
rect 38668 13022 38670 13074
rect 38722 13022 38724 13074
rect 38668 13010 38724 13022
rect 39452 12852 39508 12862
rect 39452 12758 39508 12796
rect 39676 12850 39732 12862
rect 39676 12798 39678 12850
rect 39730 12798 39732 12850
rect 39676 12404 39732 12798
rect 40236 12852 40292 12862
rect 40236 12758 40292 12796
rect 39676 12338 39732 12348
rect 37772 11172 37828 11182
rect 37772 11170 38388 11172
rect 37772 11118 37774 11170
rect 37826 11118 38388 11170
rect 37772 11116 38388 11118
rect 37772 11106 37828 11116
rect 37772 10836 37828 10846
rect 37772 10834 38276 10836
rect 37772 10782 37774 10834
rect 37826 10782 38276 10834
rect 37772 10780 38276 10782
rect 37772 10770 37828 10780
rect 35308 9538 35364 9548
rect 36204 9538 36260 9548
rect 36316 9716 36372 9726
rect 34636 9266 34916 9268
rect 34636 9214 34638 9266
rect 34690 9214 34916 9266
rect 34636 9212 34916 9214
rect 35084 9268 35140 9278
rect 34636 9202 34692 9212
rect 35084 9174 35140 9212
rect 34188 9102 34190 9154
rect 34242 9102 34244 9154
rect 34188 9090 34244 9102
rect 33964 8978 34020 8988
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 36316 8370 36372 9660
rect 36316 8318 36318 8370
rect 36370 8318 36372 8370
rect 36316 8306 36372 8318
rect 33180 8206 33182 8258
rect 33234 8206 33236 8258
rect 33180 8194 33236 8206
rect 35756 8034 35812 8046
rect 35756 7982 35758 8034
rect 35810 7982 35812 8034
rect 33180 7700 33236 7710
rect 33068 7698 33236 7700
rect 33068 7646 33182 7698
rect 33234 7646 33236 7698
rect 33068 7644 33236 7646
rect 33180 7634 33236 7644
rect 35756 7698 35812 7982
rect 35756 7646 35758 7698
rect 35810 7646 35812 7698
rect 35756 7634 35812 7646
rect 32396 7588 32452 7598
rect 31948 7586 32396 7588
rect 31948 7534 31950 7586
rect 32002 7534 32396 7586
rect 31948 7532 32396 7534
rect 31948 7522 32004 7532
rect 32396 7494 32452 7532
rect 35420 7588 35476 7598
rect 35420 7494 35476 7532
rect 35868 7588 35924 7598
rect 35868 7494 35924 7532
rect 37660 7588 37716 10668
rect 38220 10612 38276 10780
rect 38332 10834 38388 11116
rect 38332 10782 38334 10834
rect 38386 10782 38388 10834
rect 38332 10770 38388 10782
rect 38668 10724 38724 10734
rect 38668 10630 38724 10668
rect 39116 10724 39172 10734
rect 39116 10630 39172 10668
rect 38556 10612 38612 10622
rect 38220 10610 38612 10612
rect 38220 10558 38558 10610
rect 38610 10558 38612 10610
rect 38220 10556 38612 10558
rect 38556 10546 38612 10556
rect 37660 7522 37716 7532
rect 31388 7476 31444 7486
rect 31276 7474 31780 7476
rect 31276 7422 31390 7474
rect 31442 7422 31780 7474
rect 31276 7420 31780 7422
rect 30940 7410 30996 7420
rect 31388 7410 31444 7420
rect 31724 6804 31780 7420
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 31836 6804 31892 6814
rect 31724 6802 31892 6804
rect 31724 6750 31838 6802
rect 31890 6750 31892 6802
rect 31724 6748 31892 6750
rect 28364 6692 28420 6702
rect 28364 6598 28420 6636
rect 31724 6692 31780 6748
rect 31836 6738 31892 6748
rect 31724 6626 31780 6636
rect 27804 6514 27860 6524
rect 26796 6414 26798 6466
rect 26850 6414 26852 6466
rect 26796 6402 26852 6414
rect 27916 6468 27972 6478
rect 27916 6374 27972 6412
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 26908 3668 26964 3678
rect 26460 3502 26462 3554
rect 26514 3502 26516 3554
rect 26460 3490 26516 3502
rect 26572 3666 26964 3668
rect 26572 3614 26910 3666
rect 26962 3614 26964 3666
rect 26572 3612 26964 3614
rect 26012 3332 26180 3388
rect 22876 800 22932 3332
rect 26012 2548 26068 3332
rect 25564 2492 26068 2548
rect 25564 800 25620 2492
rect 26572 980 26628 3612
rect 26908 3602 26964 3612
rect 26236 924 26628 980
rect 26236 800 26292 924
rect 17164 700 17668 756
rect 18144 0 18256 800
rect 21504 0 21616 800
rect 22848 0 22960 800
rect 25536 0 25648 800
rect 26208 0 26320 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 7532 36428 7588 36484
rect 4060 36316 4116 36372
rect 3948 33852 4004 33908
rect 2044 31666 2100 31668
rect 2044 31614 2046 31666
rect 2046 31614 2098 31666
rect 2098 31614 2100 31666
rect 2044 31612 2100 31614
rect 1708 31554 1764 31556
rect 1708 31502 1710 31554
rect 1710 31502 1762 31554
rect 1762 31502 1764 31554
rect 1708 31500 1764 31502
rect 2492 31554 2548 31556
rect 2492 31502 2494 31554
rect 2494 31502 2546 31554
rect 2546 31502 2548 31554
rect 2492 31500 2548 31502
rect 3276 31500 3332 31556
rect 1708 30940 1764 30996
rect 2828 31052 2884 31108
rect 2156 30210 2212 30212
rect 2156 30158 2158 30210
rect 2158 30158 2210 30210
rect 2210 30158 2212 30210
rect 2156 30156 2212 30158
rect 1708 28924 1764 28980
rect 2492 28924 2548 28980
rect 2044 28812 2100 28868
rect 2940 28700 2996 28756
rect 2156 28418 2212 28420
rect 2156 28366 2158 28418
rect 2158 28366 2210 28418
rect 2210 28366 2212 28418
rect 2156 28364 2212 28366
rect 3836 27858 3892 27860
rect 3836 27806 3838 27858
rect 3838 27806 3890 27858
rect 3890 27806 3892 27858
rect 3836 27804 3892 27806
rect 1932 25564 1988 25620
rect 2044 25004 2100 25060
rect 2156 24892 2212 24948
rect 2940 25564 2996 25620
rect 2828 25228 2884 25284
rect 3612 24946 3668 24948
rect 3612 24894 3614 24946
rect 3614 24894 3666 24946
rect 3666 24894 3668 24946
rect 3612 24892 3668 24894
rect 1708 24220 1764 24276
rect 2492 24220 2548 24276
rect 2268 23938 2324 23940
rect 2268 23886 2270 23938
rect 2270 23886 2322 23938
rect 2322 23886 2324 23938
rect 2268 23884 2324 23886
rect 1708 23548 1764 23604
rect 2716 23548 2772 23604
rect 2828 23324 2884 23380
rect 3388 23378 3444 23380
rect 3388 23326 3390 23378
rect 3390 23326 3442 23378
rect 3442 23326 3444 23378
rect 3388 23324 3444 23326
rect 1932 23042 1988 23044
rect 1932 22990 1934 23042
rect 1934 22990 1986 23042
rect 1986 22990 1988 23042
rect 1932 22988 1988 22990
rect 1932 22258 1988 22260
rect 1932 22206 1934 22258
rect 1934 22206 1986 22258
rect 1986 22206 1988 22258
rect 1932 22204 1988 22206
rect 1596 22092 1652 22148
rect 3276 22258 3332 22260
rect 3276 22206 3278 22258
rect 3278 22206 3330 22258
rect 3330 22206 3332 22258
rect 3276 22204 3332 22206
rect 2828 22092 2884 22148
rect 2380 21810 2436 21812
rect 2380 21758 2382 21810
rect 2382 21758 2434 21810
rect 2434 21758 2436 21810
rect 2380 21756 2436 21758
rect 3836 21644 3892 21700
rect 2156 21532 2212 21588
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 6412 33628 6468 33684
rect 4284 33404 4340 33460
rect 6188 33458 6244 33460
rect 6188 33406 6190 33458
rect 6190 33406 6242 33458
rect 6242 33406 6244 33458
rect 6188 33404 6244 33406
rect 6076 33122 6132 33124
rect 6076 33070 6078 33122
rect 6078 33070 6130 33122
rect 6130 33070 6132 33122
rect 6076 33068 6132 33070
rect 6076 32450 6132 32452
rect 6076 32398 6078 32450
rect 6078 32398 6130 32450
rect 6130 32398 6132 32450
rect 6076 32396 6132 32398
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 5964 32060 6020 32116
rect 5740 31554 5796 31556
rect 5740 31502 5742 31554
rect 5742 31502 5794 31554
rect 5794 31502 5796 31554
rect 5740 31500 5796 31502
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5180 29986 5236 29988
rect 5180 29934 5182 29986
rect 5182 29934 5234 29986
rect 5234 29934 5236 29986
rect 5180 29932 5236 29934
rect 6300 32060 6356 32116
rect 6636 33516 6692 33572
rect 7420 34354 7476 34356
rect 7420 34302 7422 34354
rect 7422 34302 7474 34354
rect 7474 34302 7476 34354
rect 7420 34300 7476 34302
rect 11004 38050 11060 38052
rect 11004 37998 11006 38050
rect 11006 37998 11058 38050
rect 11058 37998 11060 38050
rect 11004 37996 11060 37998
rect 12684 38332 12740 38388
rect 14812 38220 14868 38276
rect 15484 38274 15540 38276
rect 15484 38222 15486 38274
rect 15486 38222 15538 38274
rect 15538 38222 15540 38274
rect 15484 38220 15540 38222
rect 11676 38050 11732 38052
rect 11676 37998 11678 38050
rect 11678 37998 11730 38050
rect 11730 37998 11732 38050
rect 11676 37996 11732 37998
rect 11452 37826 11508 37828
rect 11452 37774 11454 37826
rect 11454 37774 11506 37826
rect 11506 37774 11508 37826
rect 11452 37772 11508 37774
rect 9100 36482 9156 36484
rect 9100 36430 9102 36482
rect 9102 36430 9154 36482
rect 9154 36430 9156 36482
rect 9100 36428 9156 36430
rect 9548 35868 9604 35924
rect 8540 34300 8596 34356
rect 7532 33628 7588 33684
rect 8092 34076 8148 34132
rect 6972 33570 7028 33572
rect 6972 33518 6974 33570
rect 6974 33518 7026 33570
rect 7026 33518 7028 33570
rect 6972 33516 7028 33518
rect 9100 34690 9156 34692
rect 9100 34638 9102 34690
rect 9102 34638 9154 34690
rect 9154 34638 9156 34690
rect 9100 34636 9156 34638
rect 8876 34130 8932 34132
rect 8876 34078 8878 34130
rect 8878 34078 8930 34130
rect 8930 34078 8932 34130
rect 8876 34076 8932 34078
rect 9212 34076 9268 34132
rect 7868 33346 7924 33348
rect 7868 33294 7870 33346
rect 7870 33294 7922 33346
rect 7922 33294 7924 33346
rect 7868 33292 7924 33294
rect 8876 33346 8932 33348
rect 8876 33294 8878 33346
rect 8878 33294 8930 33346
rect 8930 33294 8932 33346
rect 8876 33292 8932 33294
rect 6860 32060 6916 32116
rect 8652 33122 8708 33124
rect 8652 33070 8654 33122
rect 8654 33070 8706 33122
rect 8706 33070 8708 33122
rect 8652 33068 8708 33070
rect 9772 33516 9828 33572
rect 11228 37154 11284 37156
rect 11228 37102 11230 37154
rect 11230 37102 11282 37154
rect 11282 37102 11284 37154
rect 11228 37100 11284 37102
rect 10780 36428 10836 36484
rect 12908 37100 12964 37156
rect 12572 36764 12628 36820
rect 12124 36652 12180 36708
rect 11676 36428 11732 36484
rect 11340 35922 11396 35924
rect 11340 35870 11342 35922
rect 11342 35870 11394 35922
rect 11394 35870 11396 35922
rect 11340 35868 11396 35870
rect 11004 35698 11060 35700
rect 11004 35646 11006 35698
rect 11006 35646 11058 35698
rect 11058 35646 11060 35698
rect 11004 35644 11060 35646
rect 10108 34636 10164 34692
rect 10108 34130 10164 34132
rect 10108 34078 10110 34130
rect 10110 34078 10162 34130
rect 10162 34078 10164 34130
rect 10108 34076 10164 34078
rect 11452 35698 11508 35700
rect 11452 35646 11454 35698
rect 11454 35646 11506 35698
rect 11506 35646 11508 35698
rect 11452 35644 11508 35646
rect 11676 35196 11732 35252
rect 10332 33964 10388 34020
rect 10108 33292 10164 33348
rect 9100 32732 9156 32788
rect 8988 32620 9044 32676
rect 7196 32396 7252 32452
rect 6524 31106 6580 31108
rect 6524 31054 6526 31106
rect 6526 31054 6578 31106
rect 6578 31054 6580 31106
rect 6524 31052 6580 31054
rect 8204 31836 8260 31892
rect 7308 31666 7364 31668
rect 7308 31614 7310 31666
rect 7310 31614 7362 31666
rect 7362 31614 7364 31666
rect 7308 31612 7364 31614
rect 9548 31724 9604 31780
rect 7756 31612 7812 31668
rect 6076 30210 6132 30212
rect 6076 30158 6078 30210
rect 6078 30158 6130 30210
rect 6130 30158 6132 30210
rect 6076 30156 6132 30158
rect 6300 29932 6356 29988
rect 5628 29426 5684 29428
rect 5628 29374 5630 29426
rect 5630 29374 5682 29426
rect 5682 29374 5684 29426
rect 5628 29372 5684 29374
rect 6076 29260 6132 29316
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4284 28364 4340 28420
rect 5964 28418 6020 28420
rect 5964 28366 5966 28418
rect 5966 28366 6018 28418
rect 6018 28366 6020 28418
rect 5964 28364 6020 28366
rect 6748 30210 6804 30212
rect 6748 30158 6750 30210
rect 6750 30158 6802 30210
rect 6802 30158 6804 30210
rect 6748 30156 6804 30158
rect 6524 30098 6580 30100
rect 6524 30046 6526 30098
rect 6526 30046 6578 30098
rect 6578 30046 6580 30098
rect 6524 30044 6580 30046
rect 7420 31052 7476 31108
rect 8876 31666 8932 31668
rect 8876 31614 8878 31666
rect 8878 31614 8930 31666
rect 8930 31614 8932 31666
rect 8876 31612 8932 31614
rect 7308 30098 7364 30100
rect 7308 30046 7310 30098
rect 7310 30046 7362 30098
rect 7362 30046 7364 30098
rect 7308 30044 7364 30046
rect 6636 29484 6692 29540
rect 6636 29314 6692 29316
rect 6636 29262 6638 29314
rect 6638 29262 6690 29314
rect 6690 29262 6692 29314
rect 6636 29260 6692 29262
rect 6860 28700 6916 28756
rect 5852 28140 5908 28196
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 6748 28082 6804 28084
rect 6748 28030 6750 28082
rect 6750 28030 6802 28082
rect 6802 28030 6804 28082
rect 6748 28028 6804 28030
rect 6188 27804 6244 27860
rect 6300 26908 6356 26964
rect 5628 26124 5684 26180
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4956 24892 5012 24948
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 7308 28700 7364 28756
rect 6748 25788 6804 25844
rect 7084 27804 7140 27860
rect 7980 30940 8036 30996
rect 7644 29484 7700 29540
rect 8764 31276 8820 31332
rect 8316 30156 8372 30212
rect 8540 31106 8596 31108
rect 8540 31054 8542 31106
rect 8542 31054 8594 31106
rect 8594 31054 8596 31106
rect 8540 31052 8596 31054
rect 8652 30940 8708 30996
rect 8092 29708 8148 29764
rect 8540 29932 8596 29988
rect 7644 28700 7700 28756
rect 8316 28754 8372 28756
rect 8316 28702 8318 28754
rect 8318 28702 8370 28754
rect 8370 28702 8372 28754
rect 8316 28700 8372 28702
rect 8204 28642 8260 28644
rect 8204 28590 8206 28642
rect 8206 28590 8258 28642
rect 8258 28590 8260 28642
rect 8204 28588 8260 28590
rect 7532 28082 7588 28084
rect 7532 28030 7534 28082
rect 7534 28030 7586 28082
rect 7586 28030 7588 28082
rect 7532 28028 7588 28030
rect 8092 27580 8148 27636
rect 5404 24668 5460 24724
rect 5068 22428 5124 22484
rect 4732 21756 4788 21812
rect 4060 21532 4116 21588
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4508 20972 4564 21028
rect 1708 20860 1764 20916
rect 3724 20914 3780 20916
rect 3724 20862 3726 20914
rect 3726 20862 3778 20914
rect 3778 20862 3780 20914
rect 3724 20860 3780 20862
rect 4284 20802 4340 20804
rect 4284 20750 4286 20802
rect 4286 20750 4338 20802
rect 4338 20750 4340 20802
rect 4284 20748 4340 20750
rect 2604 20188 2660 20244
rect 2268 20076 2324 20132
rect 1932 19516 1988 19572
rect 2044 19122 2100 19124
rect 2044 19070 2046 19122
rect 2046 19070 2098 19122
rect 2098 19070 2100 19122
rect 2044 19068 2100 19070
rect 4732 20690 4788 20692
rect 4732 20638 4734 20690
rect 4734 20638 4786 20690
rect 4786 20638 4788 20690
rect 4732 20636 4788 20638
rect 3612 20188 3668 20244
rect 4172 20076 4228 20132
rect 3164 19740 3220 19796
rect 2940 19234 2996 19236
rect 2940 19182 2942 19234
rect 2942 19182 2994 19234
rect 2994 19182 2996 19234
rect 2940 19180 2996 19182
rect 2716 18508 2772 18564
rect 3164 18956 3220 19012
rect 2156 18450 2212 18452
rect 2156 18398 2158 18450
rect 2158 18398 2210 18450
rect 2210 18398 2212 18450
rect 2156 18396 2212 18398
rect 1708 17554 1764 17556
rect 1708 17502 1710 17554
rect 1710 17502 1762 17554
rect 1762 17502 1764 17554
rect 1708 17500 1764 17502
rect 2604 18284 2660 18340
rect 2268 18172 2324 18228
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 3612 19122 3668 19124
rect 3612 19070 3614 19122
rect 3614 19070 3666 19122
rect 3666 19070 3668 19122
rect 3612 19068 3668 19070
rect 4508 19292 4564 19348
rect 4172 18956 4228 19012
rect 3388 18060 3444 18116
rect 3724 18508 3780 18564
rect 4620 18284 4676 18340
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 5740 22482 5796 22484
rect 5740 22430 5742 22482
rect 5742 22430 5794 22482
rect 5794 22430 5796 22482
rect 5740 22428 5796 22430
rect 5628 22092 5684 22148
rect 5740 21756 5796 21812
rect 6636 25282 6692 25284
rect 6636 25230 6638 25282
rect 6638 25230 6690 25282
rect 6690 25230 6692 25282
rect 6636 25228 6692 25230
rect 6524 24722 6580 24724
rect 6524 24670 6526 24722
rect 6526 24670 6578 24722
rect 6578 24670 6580 24722
rect 6524 24668 6580 24670
rect 8652 28812 8708 28868
rect 8876 29538 8932 29540
rect 8876 29486 8878 29538
rect 8878 29486 8930 29538
rect 8930 29486 8932 29538
rect 8876 29484 8932 29486
rect 9212 31052 9268 31108
rect 9324 30940 9380 30996
rect 9548 31276 9604 31332
rect 9660 31052 9716 31108
rect 10108 33068 10164 33124
rect 9884 32732 9940 32788
rect 10108 32620 10164 32676
rect 9884 32562 9940 32564
rect 9884 32510 9886 32562
rect 9886 32510 9938 32562
rect 9938 32510 9940 32562
rect 9884 32508 9940 32510
rect 9884 31836 9940 31892
rect 10108 31612 10164 31668
rect 11900 36258 11956 36260
rect 11900 36206 11902 36258
rect 11902 36206 11954 36258
rect 11954 36206 11956 36258
rect 11900 36204 11956 36206
rect 13916 36764 13972 36820
rect 12908 36594 12964 36596
rect 12908 36542 12910 36594
rect 12910 36542 12962 36594
rect 12962 36542 12964 36594
rect 12908 36540 12964 36542
rect 13468 36652 13524 36708
rect 13132 36428 13188 36484
rect 12796 36258 12852 36260
rect 12796 36206 12798 36258
rect 12798 36206 12850 36258
rect 12850 36206 12852 36258
rect 12796 36204 12852 36206
rect 13580 36540 13636 36596
rect 12236 35308 12292 35364
rect 11900 34076 11956 34132
rect 10556 33570 10612 33572
rect 10556 33518 10558 33570
rect 10558 33518 10610 33570
rect 10610 33518 10612 33570
rect 10556 33516 10612 33518
rect 11116 33068 11172 33124
rect 10892 32674 10948 32676
rect 10892 32622 10894 32674
rect 10894 32622 10946 32674
rect 10946 32622 10948 32674
rect 10892 32620 10948 32622
rect 11116 32508 11172 32564
rect 9772 30322 9828 30324
rect 9772 30270 9774 30322
rect 9774 30270 9826 30322
rect 9826 30270 9828 30322
rect 9772 30268 9828 30270
rect 10220 30210 10276 30212
rect 10220 30158 10222 30210
rect 10222 30158 10274 30210
rect 10274 30158 10276 30210
rect 10220 30156 10276 30158
rect 9548 29932 9604 29988
rect 9324 29596 9380 29652
rect 10220 29708 10276 29764
rect 8764 28588 8820 28644
rect 10444 30156 10500 30212
rect 11452 33964 11508 34020
rect 12012 33964 12068 34020
rect 11676 33068 11732 33124
rect 11452 32620 11508 32676
rect 11228 30604 11284 30660
rect 11004 30156 11060 30212
rect 10444 29650 10500 29652
rect 10444 29598 10446 29650
rect 10446 29598 10498 29650
rect 10498 29598 10500 29650
rect 10444 29596 10500 29598
rect 10108 29426 10164 29428
rect 10108 29374 10110 29426
rect 10110 29374 10162 29426
rect 10162 29374 10164 29426
rect 10108 29372 10164 29374
rect 10556 29426 10612 29428
rect 10556 29374 10558 29426
rect 10558 29374 10610 29426
rect 10610 29374 10612 29426
rect 10556 29372 10612 29374
rect 9884 28812 9940 28868
rect 10220 28924 10276 28980
rect 9772 28700 9828 28756
rect 10108 28754 10164 28756
rect 10108 28702 10110 28754
rect 10110 28702 10162 28754
rect 10162 28702 10164 28754
rect 10108 28700 10164 28702
rect 9660 28028 9716 28084
rect 10556 28812 10612 28868
rect 11564 31666 11620 31668
rect 11564 31614 11566 31666
rect 11566 31614 11618 31666
rect 11618 31614 11620 31666
rect 11564 31612 11620 31614
rect 11452 30994 11508 30996
rect 11452 30942 11454 30994
rect 11454 30942 11506 30994
rect 11506 30942 11508 30994
rect 11452 30940 11508 30942
rect 11452 30268 11508 30324
rect 11340 28812 11396 28868
rect 11004 28700 11060 28756
rect 10556 28588 10612 28644
rect 10444 28140 10500 28196
rect 10332 28082 10388 28084
rect 10332 28030 10334 28082
rect 10334 28030 10386 28082
rect 10386 28030 10388 28082
rect 10332 28028 10388 28030
rect 11452 28642 11508 28644
rect 11452 28590 11454 28642
rect 11454 28590 11506 28642
rect 11506 28590 11508 28642
rect 11452 28588 11508 28590
rect 10780 28364 10836 28420
rect 9212 27244 9268 27300
rect 9884 27244 9940 27300
rect 8540 27132 8596 27188
rect 7532 26402 7588 26404
rect 7532 26350 7534 26402
rect 7534 26350 7586 26402
rect 7586 26350 7588 26402
rect 7532 26348 7588 26350
rect 6860 24668 6916 24724
rect 7084 23996 7140 24052
rect 7196 23938 7252 23940
rect 7196 23886 7198 23938
rect 7198 23886 7250 23938
rect 7250 23886 7252 23938
rect 7196 23884 7252 23886
rect 7308 23100 7364 23156
rect 6412 22316 6468 22372
rect 6188 22092 6244 22148
rect 6188 21644 6244 21700
rect 5964 20748 6020 20804
rect 5180 20130 5236 20132
rect 5180 20078 5182 20130
rect 5182 20078 5234 20130
rect 5234 20078 5236 20130
rect 5180 20076 5236 20078
rect 6524 22092 6580 22148
rect 6748 21756 6804 21812
rect 6636 21644 6692 21700
rect 6188 20802 6244 20804
rect 6188 20750 6190 20802
rect 6190 20750 6242 20802
rect 6242 20750 6244 20802
rect 6188 20748 6244 20750
rect 6524 20748 6580 20804
rect 6076 20300 6132 20356
rect 5628 20130 5684 20132
rect 5628 20078 5630 20130
rect 5630 20078 5682 20130
rect 5682 20078 5684 20130
rect 5628 20076 5684 20078
rect 6412 20300 6468 20356
rect 6636 20636 6692 20692
rect 5740 19180 5796 19236
rect 6300 19234 6356 19236
rect 6300 19182 6302 19234
rect 6302 19182 6354 19234
rect 6354 19182 6356 19234
rect 6300 19180 6356 19182
rect 6188 18674 6244 18676
rect 6188 18622 6190 18674
rect 6190 18622 6242 18674
rect 6242 18622 6244 18674
rect 6188 18620 6244 18622
rect 6524 18396 6580 18452
rect 6972 20076 7028 20132
rect 8316 26348 8372 26404
rect 7980 26290 8036 26292
rect 7980 26238 7982 26290
rect 7982 26238 8034 26290
rect 8034 26238 8036 26290
rect 7980 26236 8036 26238
rect 7868 26178 7924 26180
rect 7868 26126 7870 26178
rect 7870 26126 7922 26178
rect 7922 26126 7924 26178
rect 7868 26124 7924 26126
rect 7644 25228 7700 25284
rect 7980 25116 8036 25172
rect 9548 26348 9604 26404
rect 8764 25730 8820 25732
rect 8764 25678 8766 25730
rect 8766 25678 8818 25730
rect 8818 25678 8820 25730
rect 8764 25676 8820 25678
rect 8092 23660 8148 23716
rect 8092 23212 8148 23268
rect 7532 22482 7588 22484
rect 7532 22430 7534 22482
rect 7534 22430 7586 22482
rect 7586 22430 7588 22482
rect 7532 22428 7588 22430
rect 7196 20748 7252 20804
rect 7980 22482 8036 22484
rect 7980 22430 7982 22482
rect 7982 22430 8034 22482
rect 8034 22430 8036 22482
rect 7980 22428 8036 22430
rect 8092 21980 8148 22036
rect 9660 26290 9716 26292
rect 9660 26238 9662 26290
rect 9662 26238 9714 26290
rect 9714 26238 9716 26290
rect 9660 26236 9716 26238
rect 9548 25676 9604 25732
rect 9772 25506 9828 25508
rect 9772 25454 9774 25506
rect 9774 25454 9826 25506
rect 9826 25454 9828 25506
rect 9772 25452 9828 25454
rect 8652 25228 8708 25284
rect 8540 25116 8596 25172
rect 8428 25004 8484 25060
rect 8316 23212 8372 23268
rect 8540 24050 8596 24052
rect 8540 23998 8542 24050
rect 8542 23998 8594 24050
rect 8594 23998 8596 24050
rect 8540 23996 8596 23998
rect 9548 25004 9604 25060
rect 8988 24668 9044 24724
rect 8764 23660 8820 23716
rect 8428 22540 8484 22596
rect 8428 22204 8484 22260
rect 8652 22764 8708 22820
rect 8652 22482 8708 22484
rect 8652 22430 8654 22482
rect 8654 22430 8706 22482
rect 8706 22430 8708 22482
rect 8652 22428 8708 22430
rect 8764 22316 8820 22372
rect 8876 22146 8932 22148
rect 8876 22094 8878 22146
rect 8878 22094 8930 22146
rect 8930 22094 8932 22146
rect 8876 22092 8932 22094
rect 9436 23826 9492 23828
rect 9436 23774 9438 23826
rect 9438 23774 9490 23826
rect 9490 23774 9492 23826
rect 9436 23772 9492 23774
rect 9548 23436 9604 23492
rect 9772 23660 9828 23716
rect 9660 23266 9716 23268
rect 9660 23214 9662 23266
rect 9662 23214 9714 23266
rect 9714 23214 9716 23266
rect 9660 23212 9716 23214
rect 9548 23154 9604 23156
rect 9548 23102 9550 23154
rect 9550 23102 9602 23154
rect 9602 23102 9604 23154
rect 9548 23100 9604 23102
rect 9772 22876 9828 22932
rect 9212 22764 9268 22820
rect 10444 27298 10500 27300
rect 10444 27246 10446 27298
rect 10446 27246 10498 27298
rect 10498 27246 10500 27298
rect 10444 27244 10500 27246
rect 11452 26908 11508 26964
rect 11228 26460 11284 26516
rect 11116 26348 11172 26404
rect 11340 26348 11396 26404
rect 10108 25004 10164 25060
rect 10220 24946 10276 24948
rect 10220 24894 10222 24946
rect 10222 24894 10274 24946
rect 10274 24894 10276 24946
rect 10220 24892 10276 24894
rect 9996 24722 10052 24724
rect 9996 24670 9998 24722
rect 9998 24670 10050 24722
rect 10050 24670 10052 24722
rect 9996 24668 10052 24670
rect 9996 24444 10052 24500
rect 9324 22540 9380 22596
rect 8204 20972 8260 21028
rect 7420 20690 7476 20692
rect 7420 20638 7422 20690
rect 7422 20638 7474 20690
rect 7474 20638 7476 20690
rect 7420 20636 7476 20638
rect 7644 20300 7700 20356
rect 7644 19964 7700 20020
rect 7868 20018 7924 20020
rect 7868 19966 7870 20018
rect 7870 19966 7922 20018
rect 7922 19966 7924 20018
rect 7868 19964 7924 19966
rect 7644 19628 7700 19684
rect 8428 20636 8484 20692
rect 8316 20076 8372 20132
rect 7980 19852 8036 19908
rect 7532 19404 7588 19460
rect 6860 18620 6916 18676
rect 8428 20018 8484 20020
rect 8428 19966 8430 20018
rect 8430 19966 8482 20018
rect 8482 19966 8484 20018
rect 8428 19964 8484 19966
rect 8876 20300 8932 20356
rect 9212 20636 9268 20692
rect 9436 21980 9492 22036
rect 10444 25452 10500 25508
rect 11228 25394 11284 25396
rect 11228 25342 11230 25394
rect 11230 25342 11282 25394
rect 11282 25342 11284 25394
rect 11228 25340 11284 25342
rect 10220 23436 10276 23492
rect 10668 24780 10724 24836
rect 11340 24834 11396 24836
rect 11340 24782 11342 24834
rect 11342 24782 11394 24834
rect 11394 24782 11396 24834
rect 11340 24780 11396 24782
rect 11228 24444 11284 24500
rect 10556 23938 10612 23940
rect 10556 23886 10558 23938
rect 10558 23886 10610 23938
rect 10610 23886 10612 23938
rect 10556 23884 10612 23886
rect 11564 23884 11620 23940
rect 10444 23772 10500 23828
rect 10332 23212 10388 23268
rect 11116 23212 11172 23268
rect 12460 35026 12516 35028
rect 12460 34974 12462 35026
rect 12462 34974 12514 35026
rect 12514 34974 12516 35026
rect 12460 34972 12516 34974
rect 12684 34130 12740 34132
rect 12684 34078 12686 34130
rect 12686 34078 12738 34130
rect 12738 34078 12740 34130
rect 12684 34076 12740 34078
rect 12796 34018 12852 34020
rect 12796 33966 12798 34018
rect 12798 33966 12850 34018
rect 12850 33966 12852 34018
rect 12796 33964 12852 33966
rect 12572 32732 12628 32788
rect 12796 32620 12852 32676
rect 12124 31612 12180 31668
rect 11788 30716 11844 30772
rect 11900 30210 11956 30212
rect 11900 30158 11902 30210
rect 11902 30158 11954 30210
rect 11954 30158 11956 30210
rect 11900 30156 11956 30158
rect 12572 32060 12628 32116
rect 12124 30994 12180 30996
rect 12124 30942 12126 30994
rect 12126 30942 12178 30994
rect 12178 30942 12180 30994
rect 12124 30940 12180 30942
rect 12460 30716 12516 30772
rect 12236 30210 12292 30212
rect 12236 30158 12238 30210
rect 12238 30158 12290 30210
rect 12290 30158 12292 30210
rect 12236 30156 12292 30158
rect 12796 30828 12852 30884
rect 11900 28924 11956 28980
rect 14812 36988 14868 37044
rect 15148 36876 15204 36932
rect 15932 37772 15988 37828
rect 16716 38332 16772 38388
rect 16156 37436 16212 37492
rect 17500 38332 17556 38388
rect 18172 38274 18228 38276
rect 18172 38222 18174 38274
rect 18174 38222 18226 38274
rect 18226 38222 18228 38274
rect 18172 38220 18228 38222
rect 15260 36428 15316 36484
rect 15372 36988 15428 37044
rect 13916 35980 13972 36036
rect 13916 35532 13972 35588
rect 14476 35532 14532 35588
rect 14028 34914 14084 34916
rect 14028 34862 14030 34914
rect 14030 34862 14082 34914
rect 14082 34862 14084 34914
rect 14028 34860 14084 34862
rect 13020 34690 13076 34692
rect 13020 34638 13022 34690
rect 13022 34638 13074 34690
rect 13074 34638 13076 34690
rect 13020 34636 13076 34638
rect 13692 34636 13748 34692
rect 13692 33516 13748 33572
rect 14476 34914 14532 34916
rect 14476 34862 14478 34914
rect 14478 34862 14530 34914
rect 14530 34862 14532 34914
rect 14476 34860 14532 34862
rect 15036 35420 15092 35476
rect 15708 36988 15764 37044
rect 15708 36204 15764 36260
rect 15708 35810 15764 35812
rect 15708 35758 15710 35810
rect 15710 35758 15762 35810
rect 15762 35758 15764 35810
rect 15708 35756 15764 35758
rect 14924 35084 14980 35140
rect 14700 34860 14756 34916
rect 13916 34076 13972 34132
rect 13804 33292 13860 33348
rect 13692 33180 13748 33236
rect 13580 32786 13636 32788
rect 13580 32734 13582 32786
rect 13582 32734 13634 32786
rect 13634 32734 13636 32786
rect 13580 32732 13636 32734
rect 13692 32674 13748 32676
rect 13692 32622 13694 32674
rect 13694 32622 13746 32674
rect 13746 32622 13748 32674
rect 13692 32620 13748 32622
rect 13468 32060 13524 32116
rect 14812 34748 14868 34804
rect 14700 34690 14756 34692
rect 14700 34638 14702 34690
rect 14702 34638 14754 34690
rect 14754 34638 14756 34690
rect 14700 34636 14756 34638
rect 14476 34524 14532 34580
rect 14700 34412 14756 34468
rect 15036 34076 15092 34132
rect 15260 35420 15316 35476
rect 15260 35084 15316 35140
rect 15708 35420 15764 35476
rect 15260 34690 15316 34692
rect 15260 34638 15262 34690
rect 15262 34638 15314 34690
rect 15314 34638 15316 34690
rect 15260 34636 15316 34638
rect 14028 33740 14084 33796
rect 13916 31836 13972 31892
rect 13020 31612 13076 31668
rect 13468 31666 13524 31668
rect 13468 31614 13470 31666
rect 13470 31614 13522 31666
rect 13522 31614 13524 31666
rect 13468 31612 13524 31614
rect 13692 31164 13748 31220
rect 13468 31106 13524 31108
rect 13468 31054 13470 31106
rect 13470 31054 13522 31106
rect 13522 31054 13524 31106
rect 13468 31052 13524 31054
rect 13916 31612 13972 31668
rect 14140 32060 14196 32116
rect 14588 33740 14644 33796
rect 14700 33346 14756 33348
rect 14700 33294 14702 33346
rect 14702 33294 14754 33346
rect 14754 33294 14756 33346
rect 14700 33292 14756 33294
rect 15596 34412 15652 34468
rect 16156 36876 16212 36932
rect 15932 36092 15988 36148
rect 16492 36482 16548 36484
rect 16492 36430 16494 36482
rect 16494 36430 16546 36482
rect 16546 36430 16548 36482
rect 16492 36428 16548 36430
rect 16380 36092 16436 36148
rect 16716 36204 16772 36260
rect 16044 35196 16100 35252
rect 15820 34802 15876 34804
rect 15820 34750 15822 34802
rect 15822 34750 15874 34802
rect 15874 34750 15876 34802
rect 15820 34748 15876 34750
rect 15708 34188 15764 34244
rect 15596 34130 15652 34132
rect 15596 34078 15598 34130
rect 15598 34078 15650 34130
rect 15650 34078 15652 34130
rect 15596 34076 15652 34078
rect 14364 31612 14420 31668
rect 14028 31052 14084 31108
rect 14700 31724 14756 31780
rect 14924 31836 14980 31892
rect 14924 31164 14980 31220
rect 14812 31052 14868 31108
rect 15596 31666 15652 31668
rect 15596 31614 15598 31666
rect 15598 31614 15650 31666
rect 15650 31614 15652 31666
rect 15596 31612 15652 31614
rect 15372 31218 15428 31220
rect 15372 31166 15374 31218
rect 15374 31166 15426 31218
rect 15426 31166 15428 31218
rect 15372 31164 15428 31166
rect 15260 30828 15316 30884
rect 15484 30994 15540 30996
rect 15484 30942 15486 30994
rect 15486 30942 15538 30994
rect 15538 30942 15540 30994
rect 15484 30940 15540 30942
rect 14252 30434 14308 30436
rect 14252 30382 14254 30434
rect 14254 30382 14306 30434
rect 14306 30382 14308 30434
rect 14252 30380 14308 30382
rect 14028 30156 14084 30212
rect 14476 30210 14532 30212
rect 14476 30158 14478 30210
rect 14478 30158 14530 30210
rect 14530 30158 14532 30210
rect 14476 30156 14532 30158
rect 15484 30210 15540 30212
rect 15484 30158 15486 30210
rect 15486 30158 15538 30210
rect 15538 30158 15540 30210
rect 15484 30156 15540 30158
rect 14588 29932 14644 29988
rect 14140 29820 14196 29876
rect 12460 28642 12516 28644
rect 12460 28590 12462 28642
rect 12462 28590 12514 28642
rect 12514 28590 12516 28642
rect 12460 28588 12516 28590
rect 12348 26962 12404 26964
rect 12348 26910 12350 26962
rect 12350 26910 12402 26962
rect 12402 26910 12404 26962
rect 12348 26908 12404 26910
rect 12012 25506 12068 25508
rect 12012 25454 12014 25506
rect 12014 25454 12066 25506
rect 12066 25454 12068 25506
rect 12012 25452 12068 25454
rect 14140 28812 14196 28868
rect 15484 28754 15540 28756
rect 15484 28702 15486 28754
rect 15486 28702 15538 28754
rect 15538 28702 15540 28754
rect 15484 28700 15540 28702
rect 14364 28588 14420 28644
rect 12908 27692 12964 27748
rect 13356 27692 13412 27748
rect 12572 26850 12628 26852
rect 12572 26798 12574 26850
rect 12574 26798 12626 26850
rect 12626 26798 12628 26850
rect 12572 26796 12628 26798
rect 12908 26460 12964 26516
rect 12684 26348 12740 26404
rect 12460 25452 12516 25508
rect 12572 25618 12628 25620
rect 12572 25566 12574 25618
rect 12574 25566 12626 25618
rect 12626 25566 12628 25618
rect 12572 25564 12628 25566
rect 12124 25394 12180 25396
rect 12124 25342 12126 25394
rect 12126 25342 12178 25394
rect 12178 25342 12180 25394
rect 12124 25340 12180 25342
rect 11788 25004 11844 25060
rect 12796 25282 12852 25284
rect 12796 25230 12798 25282
rect 12798 25230 12850 25282
rect 12850 25230 12852 25282
rect 12796 25228 12852 25230
rect 13468 26796 13524 26852
rect 13692 25676 13748 25732
rect 13356 25564 13412 25620
rect 13468 25228 13524 25284
rect 13244 23996 13300 24052
rect 12012 23772 12068 23828
rect 13468 23826 13524 23828
rect 13468 23774 13470 23826
rect 13470 23774 13522 23826
rect 13522 23774 13524 23826
rect 13468 23772 13524 23774
rect 13692 23660 13748 23716
rect 11676 23436 11732 23492
rect 12124 23266 12180 23268
rect 12124 23214 12126 23266
rect 12126 23214 12178 23266
rect 12178 23214 12180 23266
rect 12124 23212 12180 23214
rect 10220 22316 10276 22372
rect 9772 21868 9828 21924
rect 11340 22876 11396 22932
rect 11228 22370 11284 22372
rect 11228 22318 11230 22370
rect 11230 22318 11282 22370
rect 11282 22318 11284 22370
rect 11228 22316 11284 22318
rect 10220 21868 10276 21924
rect 10444 22146 10500 22148
rect 10444 22094 10446 22146
rect 10446 22094 10498 22146
rect 10498 22094 10500 22146
rect 10444 22092 10500 22094
rect 10892 22146 10948 22148
rect 10892 22094 10894 22146
rect 10894 22094 10946 22146
rect 10946 22094 10948 22146
rect 10892 22092 10948 22094
rect 10444 21868 10500 21924
rect 9660 20802 9716 20804
rect 9660 20750 9662 20802
rect 9662 20750 9714 20802
rect 9714 20750 9716 20802
rect 9660 20748 9716 20750
rect 8540 19458 8596 19460
rect 8540 19406 8542 19458
rect 8542 19406 8594 19458
rect 8594 19406 8596 19458
rect 8540 19404 8596 19406
rect 10108 20748 10164 20804
rect 10220 20300 10276 20356
rect 9548 20076 9604 20132
rect 8764 19292 8820 19348
rect 8764 18956 8820 19012
rect 6972 18562 7028 18564
rect 6972 18510 6974 18562
rect 6974 18510 7026 18562
rect 7026 18510 7028 18562
rect 6972 18508 7028 18510
rect 7532 18562 7588 18564
rect 7532 18510 7534 18562
rect 7534 18510 7586 18562
rect 7586 18510 7588 18562
rect 7532 18508 7588 18510
rect 9324 19010 9380 19012
rect 9324 18958 9326 19010
rect 9326 18958 9378 19010
rect 9378 18958 9380 19010
rect 9324 18956 9380 18958
rect 10332 20242 10388 20244
rect 10332 20190 10334 20242
rect 10334 20190 10386 20242
rect 10386 20190 10388 20242
rect 10332 20188 10388 20190
rect 10444 20018 10500 20020
rect 10444 19966 10446 20018
rect 10446 19966 10498 20018
rect 10498 19966 10500 20018
rect 10444 19964 10500 19966
rect 10220 19010 10276 19012
rect 10220 18958 10222 19010
rect 10222 18958 10274 19010
rect 10274 18958 10276 19010
rect 10220 18956 10276 18958
rect 9772 18508 9828 18564
rect 10220 18732 10276 18788
rect 3724 17554 3780 17556
rect 3724 17502 3726 17554
rect 3726 17502 3778 17554
rect 3778 17502 3780 17554
rect 3724 17500 3780 17502
rect 2604 17442 2660 17444
rect 2604 17390 2606 17442
rect 2606 17390 2658 17442
rect 2658 17390 2660 17442
rect 2604 17388 2660 17390
rect 4060 17442 4116 17444
rect 4060 17390 4062 17442
rect 4062 17390 4114 17442
rect 4114 17390 4116 17442
rect 4060 17388 4116 17390
rect 5068 17388 5124 17444
rect 2940 17106 2996 17108
rect 2940 17054 2942 17106
rect 2942 17054 2994 17106
rect 2994 17054 2996 17106
rect 2940 17052 2996 17054
rect 2156 16156 2212 16212
rect 2044 15484 2100 15540
rect 2604 16828 2660 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 2940 16156 2996 16212
rect 10780 20188 10836 20244
rect 10668 19068 10724 19124
rect 8540 17612 8596 17668
rect 10892 20076 10948 20132
rect 10892 19906 10948 19908
rect 10892 19854 10894 19906
rect 10894 19854 10946 19906
rect 10946 19854 10948 19906
rect 10892 19852 10948 19854
rect 10892 19180 10948 19236
rect 11004 19068 11060 19124
rect 10780 18732 10836 18788
rect 10332 17612 10388 17668
rect 8540 17276 8596 17332
rect 7308 16716 7364 16772
rect 9100 17276 9156 17332
rect 9548 17388 9604 17444
rect 8988 16716 9044 16772
rect 9996 17052 10052 17108
rect 10108 16940 10164 16996
rect 10668 17612 10724 17668
rect 10780 18396 10836 18452
rect 10444 17052 10500 17108
rect 10780 17052 10836 17108
rect 11004 17724 11060 17780
rect 10892 16604 10948 16660
rect 11340 21868 11396 21924
rect 12908 22428 12964 22484
rect 11900 22204 11956 22260
rect 11452 21644 11508 21700
rect 12684 22370 12740 22372
rect 12684 22318 12686 22370
rect 12686 22318 12738 22370
rect 12738 22318 12740 22370
rect 12684 22316 12740 22318
rect 12572 21698 12628 21700
rect 12572 21646 12574 21698
rect 12574 21646 12626 21698
rect 12626 21646 12628 21698
rect 12572 21644 12628 21646
rect 13692 22428 13748 22484
rect 13468 22092 13524 22148
rect 12908 21810 12964 21812
rect 12908 21758 12910 21810
rect 12910 21758 12962 21810
rect 12962 21758 12964 21810
rect 12908 21756 12964 21758
rect 15148 28642 15204 28644
rect 15148 28590 15150 28642
rect 15150 28590 15202 28642
rect 15202 28590 15204 28642
rect 15148 28588 15204 28590
rect 16492 35698 16548 35700
rect 16492 35646 16494 35698
rect 16494 35646 16546 35698
rect 16546 35646 16548 35698
rect 16492 35644 16548 35646
rect 16492 35308 16548 35364
rect 16380 35196 16436 35252
rect 16380 34972 16436 35028
rect 16044 34914 16100 34916
rect 16044 34862 16046 34914
rect 16046 34862 16098 34914
rect 16098 34862 16100 34914
rect 16044 34860 16100 34862
rect 16268 34748 16324 34804
rect 16492 34914 16548 34916
rect 16492 34862 16494 34914
rect 16494 34862 16546 34914
rect 16546 34862 16548 34914
rect 16492 34860 16548 34862
rect 17388 37490 17444 37492
rect 17388 37438 17390 37490
rect 17390 37438 17442 37490
rect 17442 37438 17444 37490
rect 17388 37436 17444 37438
rect 16828 35644 16884 35700
rect 17836 35698 17892 35700
rect 17836 35646 17838 35698
rect 17838 35646 17890 35698
rect 17890 35646 17892 35698
rect 17836 35644 17892 35646
rect 17164 35420 17220 35476
rect 16828 34914 16884 34916
rect 16828 34862 16830 34914
rect 16830 34862 16882 34914
rect 16882 34862 16884 34914
rect 16828 34860 16884 34862
rect 16380 34636 16436 34692
rect 16940 34354 16996 34356
rect 16940 34302 16942 34354
rect 16942 34302 16994 34354
rect 16994 34302 16996 34354
rect 16940 34300 16996 34302
rect 16604 33964 16660 34020
rect 16604 33516 16660 33572
rect 16604 33346 16660 33348
rect 16604 33294 16606 33346
rect 16606 33294 16658 33346
rect 16658 33294 16660 33346
rect 16604 33292 16660 33294
rect 17052 33404 17108 33460
rect 16716 33180 16772 33236
rect 16156 30098 16212 30100
rect 16156 30046 16158 30098
rect 16158 30046 16210 30098
rect 16210 30046 16212 30098
rect 16156 30044 16212 30046
rect 16156 29426 16212 29428
rect 16156 29374 16158 29426
rect 16158 29374 16210 29426
rect 16210 29374 16212 29426
rect 16156 29372 16212 29374
rect 17388 35586 17444 35588
rect 17388 35534 17390 35586
rect 17390 35534 17442 35586
rect 17442 35534 17444 35586
rect 17388 35532 17444 35534
rect 18060 36092 18116 36148
rect 17948 35532 18004 35588
rect 19516 38220 19572 38276
rect 18620 36316 18676 36372
rect 18620 35980 18676 36036
rect 18284 35868 18340 35924
rect 17500 34914 17556 34916
rect 17500 34862 17502 34914
rect 17502 34862 17554 34914
rect 17554 34862 17556 34914
rect 17500 34860 17556 34862
rect 17388 34188 17444 34244
rect 18172 34860 18228 34916
rect 18284 35644 18340 35700
rect 18396 35084 18452 35140
rect 18844 34972 18900 35028
rect 18732 34860 18788 34916
rect 18620 34690 18676 34692
rect 18620 34638 18622 34690
rect 18622 34638 18674 34690
rect 18674 34638 18676 34690
rect 18620 34636 18676 34638
rect 17724 34300 17780 34356
rect 17836 33516 17892 33572
rect 18508 34354 18564 34356
rect 18508 34302 18510 34354
rect 18510 34302 18562 34354
rect 18562 34302 18564 34354
rect 18508 34300 18564 34302
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19180 35868 19236 35924
rect 19516 37266 19572 37268
rect 19516 37214 19518 37266
rect 19518 37214 19570 37266
rect 19570 37214 19572 37266
rect 19516 37212 19572 37214
rect 20524 36370 20580 36372
rect 20524 36318 20526 36370
rect 20526 36318 20578 36370
rect 20578 36318 20580 36370
rect 20524 36316 20580 36318
rect 19628 36258 19684 36260
rect 19628 36206 19630 36258
rect 19630 36206 19682 36258
rect 19682 36206 19684 36258
rect 19628 36204 19684 36206
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19180 35084 19236 35140
rect 18844 34188 18900 34244
rect 18396 33234 18452 33236
rect 18396 33182 18398 33234
rect 18398 33182 18450 33234
rect 18450 33182 18452 33234
rect 18396 33180 18452 33182
rect 17836 32508 17892 32564
rect 16828 31612 16884 31668
rect 16716 31218 16772 31220
rect 16716 31166 16718 31218
rect 16718 31166 16770 31218
rect 16770 31166 16772 31218
rect 16716 31164 16772 31166
rect 16604 30828 16660 30884
rect 17276 31778 17332 31780
rect 17276 31726 17278 31778
rect 17278 31726 17330 31778
rect 17330 31726 17332 31778
rect 17276 31724 17332 31726
rect 16380 29596 16436 29652
rect 16268 29260 16324 29316
rect 16716 28866 16772 28868
rect 16716 28814 16718 28866
rect 16718 28814 16770 28866
rect 16770 28814 16772 28866
rect 16716 28812 16772 28814
rect 16828 29372 16884 29428
rect 16828 28700 16884 28756
rect 16268 28530 16324 28532
rect 16268 28478 16270 28530
rect 16270 28478 16322 28530
rect 16322 28478 16324 28530
rect 16268 28476 16324 28478
rect 15932 28028 15988 28084
rect 16604 28082 16660 28084
rect 16604 28030 16606 28082
rect 16606 28030 16658 28082
rect 16658 28030 16660 28082
rect 16604 28028 16660 28030
rect 15932 27746 15988 27748
rect 15932 27694 15934 27746
rect 15934 27694 15986 27746
rect 15986 27694 15988 27746
rect 15932 27692 15988 27694
rect 14812 27580 14868 27636
rect 15260 26236 15316 26292
rect 14924 25564 14980 25620
rect 15372 25564 15428 25620
rect 15932 26290 15988 26292
rect 15932 26238 15934 26290
rect 15934 26238 15986 26290
rect 15986 26238 15988 26290
rect 15932 26236 15988 26238
rect 15820 25676 15876 25732
rect 15708 25282 15764 25284
rect 15708 25230 15710 25282
rect 15710 25230 15762 25282
rect 15762 25230 15764 25282
rect 15708 25228 15764 25230
rect 16940 30044 16996 30100
rect 18396 32620 18452 32676
rect 18844 33068 18900 33124
rect 18396 31666 18452 31668
rect 18396 31614 18398 31666
rect 18398 31614 18450 31666
rect 18450 31614 18452 31666
rect 18396 31612 18452 31614
rect 18284 31164 18340 31220
rect 18508 31106 18564 31108
rect 18508 31054 18510 31106
rect 18510 31054 18562 31106
rect 18562 31054 18564 31106
rect 18508 31052 18564 31054
rect 17500 30994 17556 30996
rect 17500 30942 17502 30994
rect 17502 30942 17554 30994
rect 17554 30942 17556 30994
rect 17500 30940 17556 30942
rect 17052 29820 17108 29876
rect 17164 30828 17220 30884
rect 17388 30322 17444 30324
rect 17388 30270 17390 30322
rect 17390 30270 17442 30322
rect 17442 30270 17444 30322
rect 17388 30268 17444 30270
rect 17164 30210 17220 30212
rect 17164 30158 17166 30210
rect 17166 30158 17218 30210
rect 17218 30158 17220 30210
rect 17164 30156 17220 30158
rect 18060 30828 18116 30884
rect 17724 30044 17780 30100
rect 17612 29820 17668 29876
rect 17164 29596 17220 29652
rect 17388 29372 17444 29428
rect 17612 29372 17668 29428
rect 17724 28812 17780 28868
rect 17276 28530 17332 28532
rect 17276 28478 17278 28530
rect 17278 28478 17330 28530
rect 17330 28478 17332 28530
rect 17276 28476 17332 28478
rect 17164 28418 17220 28420
rect 17164 28366 17166 28418
rect 17166 28366 17218 28418
rect 17218 28366 17220 28418
rect 17164 28364 17220 28366
rect 16940 26908 16996 26964
rect 16492 26290 16548 26292
rect 16492 26238 16494 26290
rect 16494 26238 16546 26290
rect 16546 26238 16548 26290
rect 16492 26236 16548 26238
rect 15820 25116 15876 25172
rect 14476 24050 14532 24052
rect 14476 23998 14478 24050
rect 14478 23998 14530 24050
rect 14530 23998 14532 24050
rect 14476 23996 14532 23998
rect 13468 21308 13524 21364
rect 11676 18732 11732 18788
rect 11452 18396 11508 18452
rect 11340 18172 11396 18228
rect 11452 17948 11508 18004
rect 11452 17778 11508 17780
rect 11452 17726 11454 17778
rect 11454 17726 11506 17778
rect 11506 17726 11508 17778
rect 11452 17724 11508 17726
rect 12348 20802 12404 20804
rect 12348 20750 12350 20802
rect 12350 20750 12402 20802
rect 12402 20750 12404 20802
rect 12348 20748 12404 20750
rect 13468 20802 13524 20804
rect 13468 20750 13470 20802
rect 13470 20750 13522 20802
rect 13522 20750 13524 20802
rect 13468 20748 13524 20750
rect 16380 24668 16436 24724
rect 15148 23660 15204 23716
rect 14028 21756 14084 21812
rect 14700 22092 14756 22148
rect 12236 19628 12292 19684
rect 12012 18396 12068 18452
rect 12460 19292 12516 19348
rect 12908 19234 12964 19236
rect 12908 19182 12910 19234
rect 12910 19182 12962 19234
rect 12962 19182 12964 19234
rect 12908 19180 12964 19182
rect 12684 19068 12740 19124
rect 12796 18396 12852 18452
rect 12572 18338 12628 18340
rect 12572 18286 12574 18338
rect 12574 18286 12626 18338
rect 12626 18286 12628 18338
rect 12572 18284 12628 18286
rect 12236 18060 12292 18116
rect 11788 17666 11844 17668
rect 11788 17614 11790 17666
rect 11790 17614 11842 17666
rect 11842 17614 11844 17666
rect 11788 17612 11844 17614
rect 12012 17276 12068 17332
rect 11900 17052 11956 17108
rect 11228 16492 11284 16548
rect 11116 15932 11172 15988
rect 9548 15484 9604 15540
rect 10108 15538 10164 15540
rect 10108 15486 10110 15538
rect 10110 15486 10162 15538
rect 10162 15486 10164 15538
rect 10108 15484 10164 15486
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 10108 14476 10164 14532
rect 7532 14418 7588 14420
rect 7532 14366 7534 14418
rect 7534 14366 7586 14418
rect 7586 14366 7588 14418
rect 7532 14364 7588 14366
rect 8428 14418 8484 14420
rect 8428 14366 8430 14418
rect 8430 14366 8482 14418
rect 8482 14366 8484 14418
rect 8428 14364 8484 14366
rect 7196 14252 7252 14308
rect 2940 13804 2996 13860
rect 5068 13858 5124 13860
rect 5068 13806 5070 13858
rect 5070 13806 5122 13858
rect 5122 13806 5124 13858
rect 5068 13804 5124 13806
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 5068 13132 5124 13188
rect 6076 13634 6132 13636
rect 6076 13582 6078 13634
rect 6078 13582 6130 13634
rect 6130 13582 6132 13634
rect 6076 13580 6132 13582
rect 7196 13580 7252 13636
rect 6524 13132 6580 13188
rect 7868 14306 7924 14308
rect 7868 14254 7870 14306
rect 7870 14254 7922 14306
rect 7922 14254 7924 14306
rect 7868 14252 7924 14254
rect 8988 13746 9044 13748
rect 8988 13694 8990 13746
rect 8990 13694 9042 13746
rect 9042 13694 9044 13746
rect 8988 13692 9044 13694
rect 9660 13692 9716 13748
rect 12460 16882 12516 16884
rect 12460 16830 12462 16882
rect 12462 16830 12514 16882
rect 12514 16830 12516 16882
rect 12460 16828 12516 16830
rect 12460 16604 12516 16660
rect 12908 18844 12964 18900
rect 12684 17500 12740 17556
rect 14924 21362 14980 21364
rect 14924 21310 14926 21362
rect 14926 21310 14978 21362
rect 14978 21310 14980 21362
rect 14924 21308 14980 21310
rect 14252 20636 14308 20692
rect 14028 20242 14084 20244
rect 14028 20190 14030 20242
rect 14030 20190 14082 20242
rect 14082 20190 14084 20242
rect 14028 20188 14084 20190
rect 14476 21026 14532 21028
rect 14476 20974 14478 21026
rect 14478 20974 14530 21026
rect 14530 20974 14532 21026
rect 14476 20972 14532 20974
rect 13916 19292 13972 19348
rect 13468 19180 13524 19236
rect 13356 18732 13412 18788
rect 12796 18060 12852 18116
rect 12572 16268 12628 16324
rect 11900 15932 11956 15988
rect 13020 17836 13076 17892
rect 13916 19122 13972 19124
rect 13916 19070 13918 19122
rect 13918 19070 13970 19122
rect 13970 19070 13972 19122
rect 13916 19068 13972 19070
rect 13692 18844 13748 18900
rect 14028 18732 14084 18788
rect 13468 17948 13524 18004
rect 13468 17724 13524 17780
rect 13468 17500 13524 17556
rect 14252 19740 14308 19796
rect 14588 19964 14644 20020
rect 14588 19068 14644 19124
rect 14700 18844 14756 18900
rect 15036 19740 15092 19796
rect 16380 23548 16436 23604
rect 16828 24610 16884 24612
rect 16828 24558 16830 24610
rect 16830 24558 16882 24610
rect 16882 24558 16884 24610
rect 16828 24556 16884 24558
rect 15372 23100 15428 23156
rect 16828 23324 16884 23380
rect 16268 22930 16324 22932
rect 16268 22878 16270 22930
rect 16270 22878 16322 22930
rect 16322 22878 16324 22930
rect 16268 22876 16324 22878
rect 15932 22428 15988 22484
rect 16604 22258 16660 22260
rect 16604 22206 16606 22258
rect 16606 22206 16658 22258
rect 16658 22206 16660 22258
rect 16604 22204 16660 22206
rect 16492 21644 16548 21700
rect 16828 21644 16884 21700
rect 15932 20972 15988 21028
rect 15708 20860 15764 20916
rect 15820 20076 15876 20132
rect 16044 20524 16100 20580
rect 15148 19404 15204 19460
rect 15036 19292 15092 19348
rect 15372 19292 15428 19348
rect 15260 18450 15316 18452
rect 15260 18398 15262 18450
rect 15262 18398 15314 18450
rect 15314 18398 15316 18450
rect 15260 18396 15316 18398
rect 14364 18172 14420 18228
rect 14252 17836 14308 17892
rect 14140 17778 14196 17780
rect 14140 17726 14142 17778
rect 14142 17726 14194 17778
rect 14194 17726 14196 17778
rect 14140 17724 14196 17726
rect 14364 17554 14420 17556
rect 14364 17502 14366 17554
rect 14366 17502 14418 17554
rect 14418 17502 14420 17554
rect 14364 17500 14420 17502
rect 14700 17724 14756 17780
rect 14028 17388 14084 17444
rect 13244 17052 13300 17108
rect 13468 16322 13524 16324
rect 13468 16270 13470 16322
rect 13470 16270 13522 16322
rect 13522 16270 13524 16322
rect 13468 16268 13524 16270
rect 13916 16882 13972 16884
rect 13916 16830 13918 16882
rect 13918 16830 13970 16882
rect 13970 16830 13972 16882
rect 13916 16828 13972 16830
rect 13580 16210 13636 16212
rect 13580 16158 13582 16210
rect 13582 16158 13634 16210
rect 13634 16158 13636 16210
rect 13580 16156 13636 16158
rect 13580 15538 13636 15540
rect 13580 15486 13582 15538
rect 13582 15486 13634 15538
rect 13634 15486 13636 15538
rect 13580 15484 13636 15486
rect 14252 16994 14308 16996
rect 14252 16942 14254 16994
rect 14254 16942 14306 16994
rect 14306 16942 14308 16994
rect 14252 16940 14308 16942
rect 15372 17612 15428 17668
rect 14924 17554 14980 17556
rect 14924 17502 14926 17554
rect 14926 17502 14978 17554
rect 14978 17502 14980 17554
rect 14924 17500 14980 17502
rect 15372 17442 15428 17444
rect 15372 17390 15374 17442
rect 15374 17390 15426 17442
rect 15426 17390 15428 17442
rect 15372 17388 15428 17390
rect 15820 19404 15876 19460
rect 16044 19292 16100 19348
rect 16380 20412 16436 20468
rect 16716 19964 16772 20020
rect 18172 30994 18228 30996
rect 18172 30942 18174 30994
rect 18174 30942 18226 30994
rect 18226 30942 18228 30994
rect 18172 30940 18228 30942
rect 18732 31554 18788 31556
rect 18732 31502 18734 31554
rect 18734 31502 18786 31554
rect 18786 31502 18788 31554
rect 18732 31500 18788 31502
rect 18732 30828 18788 30884
rect 19180 34188 19236 34244
rect 19628 35810 19684 35812
rect 19628 35758 19630 35810
rect 19630 35758 19682 35810
rect 19682 35758 19684 35810
rect 19628 35756 19684 35758
rect 20412 36258 20468 36260
rect 20412 36206 20414 36258
rect 20414 36206 20466 36258
rect 20466 36206 20468 36258
rect 20412 36204 20468 36206
rect 20972 36204 21028 36260
rect 20412 35980 20468 36036
rect 19740 35698 19796 35700
rect 19740 35646 19742 35698
rect 19742 35646 19794 35698
rect 19794 35646 19796 35698
rect 19740 35644 19796 35646
rect 20300 35644 20356 35700
rect 19852 35308 19908 35364
rect 20748 35586 20804 35588
rect 20748 35534 20750 35586
rect 20750 35534 20802 35586
rect 20802 35534 20804 35586
rect 20748 35532 20804 35534
rect 21532 36258 21588 36260
rect 21532 36206 21534 36258
rect 21534 36206 21586 36258
rect 21586 36206 21588 36258
rect 21532 36204 21588 36206
rect 21532 35980 21588 36036
rect 21756 36316 21812 36372
rect 20972 35308 21028 35364
rect 20748 35138 20804 35140
rect 20748 35086 20750 35138
rect 20750 35086 20802 35138
rect 20802 35086 20804 35138
rect 20748 35084 20804 35086
rect 20636 35026 20692 35028
rect 20636 34974 20638 35026
rect 20638 34974 20690 35026
rect 20690 34974 20692 35026
rect 20636 34972 20692 34974
rect 20300 34748 20356 34804
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19068 33458 19124 33460
rect 19068 33406 19070 33458
rect 19070 33406 19122 33458
rect 19122 33406 19124 33458
rect 19068 33404 19124 33406
rect 19180 33122 19236 33124
rect 19180 33070 19182 33122
rect 19182 33070 19234 33122
rect 19234 33070 19236 33122
rect 19180 33068 19236 33070
rect 19404 33122 19460 33124
rect 19404 33070 19406 33122
rect 19406 33070 19458 33122
rect 19458 33070 19460 33122
rect 19404 33068 19460 33070
rect 19292 32674 19348 32676
rect 19292 32622 19294 32674
rect 19294 32622 19346 32674
rect 19346 32622 19348 32674
rect 19292 32620 19348 32622
rect 19404 32562 19460 32564
rect 19404 32510 19406 32562
rect 19406 32510 19458 32562
rect 19458 32510 19460 32562
rect 19404 32508 19460 32510
rect 18956 30994 19012 30996
rect 18956 30942 18958 30994
rect 18958 30942 19010 30994
rect 19010 30942 19012 30994
rect 18956 30940 19012 30942
rect 20972 34860 21028 34916
rect 21308 35698 21364 35700
rect 21308 35646 21310 35698
rect 21310 35646 21362 35698
rect 21362 35646 21364 35698
rect 21308 35644 21364 35646
rect 21308 35308 21364 35364
rect 19964 33122 20020 33124
rect 19964 33070 19966 33122
rect 19966 33070 20018 33122
rect 20018 33070 20020 33122
rect 19964 33068 20020 33070
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20188 32396 20244 32452
rect 19516 31724 19572 31780
rect 18508 30268 18564 30324
rect 18620 30380 18676 30436
rect 18284 30156 18340 30212
rect 17948 29596 18004 29652
rect 18172 30044 18228 30100
rect 18732 30156 18788 30212
rect 17948 28754 18004 28756
rect 17948 28702 17950 28754
rect 17950 28702 18002 28754
rect 18002 28702 18004 28754
rect 17948 28700 18004 28702
rect 18620 28700 18676 28756
rect 18396 28418 18452 28420
rect 18396 28366 18398 28418
rect 18398 28366 18450 28418
rect 18450 28366 18452 28418
rect 18396 28364 18452 28366
rect 17388 26962 17444 26964
rect 17388 26910 17390 26962
rect 17390 26910 17442 26962
rect 17442 26910 17444 26962
rect 17388 26908 17444 26910
rect 18284 28028 18340 28084
rect 18396 27132 18452 27188
rect 17724 26460 17780 26516
rect 17948 26796 18004 26852
rect 17052 25452 17108 25508
rect 17276 24892 17332 24948
rect 17388 24722 17444 24724
rect 17388 24670 17390 24722
rect 17390 24670 17442 24722
rect 17442 24670 17444 24722
rect 17388 24668 17444 24670
rect 17500 24556 17556 24612
rect 18060 25004 18116 25060
rect 17276 23548 17332 23604
rect 18060 23772 18116 23828
rect 17500 23266 17556 23268
rect 17500 23214 17502 23266
rect 17502 23214 17554 23266
rect 17554 23214 17556 23266
rect 17500 23212 17556 23214
rect 17164 22258 17220 22260
rect 17164 22206 17166 22258
rect 17166 22206 17218 22258
rect 17218 22206 17220 22258
rect 17164 22204 17220 22206
rect 17052 21420 17108 21476
rect 17052 20802 17108 20804
rect 17052 20750 17054 20802
rect 17054 20750 17106 20802
rect 17106 20750 17108 20802
rect 17052 20748 17108 20750
rect 17724 23100 17780 23156
rect 17388 22146 17444 22148
rect 17388 22094 17390 22146
rect 17390 22094 17442 22146
rect 17442 22094 17444 22146
rect 17388 22092 17444 22094
rect 17500 21810 17556 21812
rect 17500 21758 17502 21810
rect 17502 21758 17554 21810
rect 17554 21758 17556 21810
rect 17500 21756 17556 21758
rect 18060 22876 18116 22932
rect 18172 22146 18228 22148
rect 18172 22094 18174 22146
rect 18174 22094 18226 22146
rect 18226 22094 18228 22146
rect 18172 22092 18228 22094
rect 17724 21756 17780 21812
rect 17948 21980 18004 22036
rect 18732 27132 18788 27188
rect 19180 30380 19236 30436
rect 19292 31666 19348 31668
rect 19292 31614 19294 31666
rect 19294 31614 19346 31666
rect 19346 31614 19348 31666
rect 19292 31612 19348 31614
rect 19740 31612 19796 31668
rect 19516 31500 19572 31556
rect 19516 31218 19572 31220
rect 19516 31166 19518 31218
rect 19518 31166 19570 31218
rect 19570 31166 19572 31218
rect 19516 31164 19572 31166
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20972 32450 21028 32452
rect 20972 32398 20974 32450
rect 20974 32398 21026 32450
rect 21026 32398 21028 32450
rect 20972 32396 21028 32398
rect 20524 31724 20580 31780
rect 19404 29932 19460 29988
rect 19292 29596 19348 29652
rect 20748 31724 20804 31780
rect 20636 31164 20692 31220
rect 20076 30210 20132 30212
rect 20076 30158 20078 30210
rect 20078 30158 20130 30210
rect 20130 30158 20132 30210
rect 20076 30156 20132 30158
rect 19516 29708 19572 29764
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19068 29538 19124 29540
rect 19068 29486 19070 29538
rect 19070 29486 19122 29538
rect 19122 29486 19124 29538
rect 19068 29484 19124 29486
rect 20300 29986 20356 29988
rect 20300 29934 20302 29986
rect 20302 29934 20354 29986
rect 20354 29934 20356 29986
rect 20300 29932 20356 29934
rect 20524 29932 20580 29988
rect 20412 29650 20468 29652
rect 20412 29598 20414 29650
rect 20414 29598 20466 29650
rect 20466 29598 20468 29650
rect 20412 29596 20468 29598
rect 20188 29484 20244 29540
rect 19180 28364 19236 28420
rect 19068 27858 19124 27860
rect 19068 27806 19070 27858
rect 19070 27806 19122 27858
rect 19122 27806 19124 27858
rect 19068 27804 19124 27806
rect 19068 27020 19124 27076
rect 19964 29372 20020 29428
rect 21308 30434 21364 30436
rect 21308 30382 21310 30434
rect 21310 30382 21362 30434
rect 21362 30382 21364 30434
rect 21308 30380 21364 30382
rect 21756 35698 21812 35700
rect 21756 35646 21758 35698
rect 21758 35646 21810 35698
rect 21810 35646 21812 35698
rect 21756 35644 21812 35646
rect 22204 37548 22260 37604
rect 22092 35980 22148 36036
rect 21980 34972 22036 35028
rect 21756 34860 21812 34916
rect 22316 35532 22372 35588
rect 22428 34972 22484 35028
rect 22428 34412 22484 34468
rect 22092 33964 22148 34020
rect 21868 33234 21924 33236
rect 21868 33182 21870 33234
rect 21870 33182 21922 33234
rect 21922 33182 21924 33234
rect 21868 33180 21924 33182
rect 21980 33068 22036 33124
rect 21868 32396 21924 32452
rect 20300 29426 20356 29428
rect 20300 29374 20302 29426
rect 20302 29374 20354 29426
rect 20354 29374 20356 29426
rect 20300 29372 20356 29374
rect 20972 29932 21028 29988
rect 20972 29314 21028 29316
rect 20972 29262 20974 29314
rect 20974 29262 21026 29314
rect 21026 29262 21028 29314
rect 20972 29260 21028 29262
rect 19964 28754 20020 28756
rect 19964 28702 19966 28754
rect 19966 28702 20018 28754
rect 20018 28702 20020 28754
rect 19964 28700 20020 28702
rect 22316 34130 22372 34132
rect 22316 34078 22318 34130
rect 22318 34078 22370 34130
rect 22370 34078 22372 34130
rect 22316 34076 22372 34078
rect 22204 32396 22260 32452
rect 22428 32172 22484 32228
rect 21980 31948 22036 32004
rect 22428 31778 22484 31780
rect 22428 31726 22430 31778
rect 22430 31726 22482 31778
rect 22482 31726 22484 31778
rect 22428 31724 22484 31726
rect 22204 31612 22260 31668
rect 22092 30156 22148 30212
rect 22988 36370 23044 36372
rect 22988 36318 22990 36370
rect 22990 36318 23042 36370
rect 23042 36318 23044 36370
rect 22988 36316 23044 36318
rect 23548 37212 23604 37268
rect 22652 35084 22708 35140
rect 26236 38556 26292 38612
rect 23660 36764 23716 36820
rect 23996 37548 24052 37604
rect 23884 36316 23940 36372
rect 25228 37378 25284 37380
rect 25228 37326 25230 37378
rect 25230 37326 25282 37378
rect 25282 37326 25284 37378
rect 25228 37324 25284 37326
rect 24668 36764 24724 36820
rect 25340 36988 25396 37044
rect 24220 36482 24276 36484
rect 24220 36430 24222 36482
rect 24222 36430 24274 36482
rect 24274 36430 24276 36482
rect 24220 36428 24276 36430
rect 22988 35026 23044 35028
rect 22988 34974 22990 35026
rect 22990 34974 23042 35026
rect 23042 34974 23044 35026
rect 22988 34972 23044 34974
rect 23436 34914 23492 34916
rect 23436 34862 23438 34914
rect 23438 34862 23490 34914
rect 23490 34862 23492 34914
rect 23436 34860 23492 34862
rect 23436 34412 23492 34468
rect 22764 34188 22820 34244
rect 23324 34300 23380 34356
rect 22652 34076 22708 34132
rect 25340 36428 25396 36484
rect 25788 37324 25844 37380
rect 24220 35698 24276 35700
rect 24220 35646 24222 35698
rect 24222 35646 24274 35698
rect 24274 35646 24276 35698
rect 24220 35644 24276 35646
rect 24220 34914 24276 34916
rect 24220 34862 24222 34914
rect 24222 34862 24274 34914
rect 24274 34862 24276 34914
rect 24220 34860 24276 34862
rect 24332 35196 24388 35252
rect 24556 35026 24612 35028
rect 24556 34974 24558 35026
rect 24558 34974 24610 35026
rect 24610 34974 24612 35026
rect 24556 34972 24612 34974
rect 24556 34802 24612 34804
rect 24556 34750 24558 34802
rect 24558 34750 24610 34802
rect 24610 34750 24612 34802
rect 24556 34748 24612 34750
rect 23660 34300 23716 34356
rect 24108 34130 24164 34132
rect 24108 34078 24110 34130
rect 24110 34078 24162 34130
rect 24162 34078 24164 34130
rect 24108 34076 24164 34078
rect 23996 33852 24052 33908
rect 24332 33964 24388 34020
rect 24780 34412 24836 34468
rect 24668 34130 24724 34132
rect 24668 34078 24670 34130
rect 24670 34078 24722 34130
rect 24722 34078 24724 34130
rect 24668 34076 24724 34078
rect 24892 34076 24948 34132
rect 23996 33346 24052 33348
rect 23996 33294 23998 33346
rect 23998 33294 24050 33346
rect 24050 33294 24052 33346
rect 23996 33292 24052 33294
rect 24220 33180 24276 33236
rect 25228 34972 25284 35028
rect 25228 34802 25284 34804
rect 25228 34750 25230 34802
rect 25230 34750 25282 34802
rect 25282 34750 25284 34802
rect 25228 34748 25284 34750
rect 25116 34300 25172 34356
rect 25228 34130 25284 34132
rect 25228 34078 25230 34130
rect 25230 34078 25282 34130
rect 25282 34078 25284 34130
rect 25228 34076 25284 34078
rect 24108 32674 24164 32676
rect 24108 32622 24110 32674
rect 24110 32622 24162 32674
rect 24162 32622 24164 32674
rect 24108 32620 24164 32622
rect 22764 32172 22820 32228
rect 22652 31948 22708 32004
rect 22204 30044 22260 30100
rect 22316 30604 22372 30660
rect 22092 29820 22148 29876
rect 21644 29596 21700 29652
rect 19628 28364 19684 28420
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 21196 27804 21252 27860
rect 19404 27074 19460 27076
rect 19404 27022 19406 27074
rect 19406 27022 19458 27074
rect 19458 27022 19460 27074
rect 19404 27020 19460 27022
rect 21980 27580 22036 27636
rect 19292 26796 19348 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 18844 25676 18900 25732
rect 18732 25116 18788 25172
rect 18732 24946 18788 24948
rect 18732 24894 18734 24946
rect 18734 24894 18786 24946
rect 18786 24894 18788 24946
rect 18732 24892 18788 24894
rect 19068 24892 19124 24948
rect 18620 24722 18676 24724
rect 18620 24670 18622 24722
rect 18622 24670 18674 24722
rect 18674 24670 18676 24722
rect 18620 24668 18676 24670
rect 18732 23826 18788 23828
rect 18732 23774 18734 23826
rect 18734 23774 18786 23826
rect 18786 23774 18788 23826
rect 18732 23772 18788 23774
rect 18620 23660 18676 23716
rect 18396 23378 18452 23380
rect 18396 23326 18398 23378
rect 18398 23326 18450 23378
rect 18450 23326 18452 23378
rect 18396 23324 18452 23326
rect 18396 23100 18452 23156
rect 17948 21644 18004 21700
rect 17612 21196 17668 21252
rect 17052 20188 17108 20244
rect 16268 18450 16324 18452
rect 16268 18398 16270 18450
rect 16270 18398 16322 18450
rect 16322 18398 16324 18450
rect 16268 18396 16324 18398
rect 16828 19234 16884 19236
rect 16828 19182 16830 19234
rect 16830 19182 16882 19234
rect 16882 19182 16884 19234
rect 16828 19180 16884 19182
rect 16492 18396 16548 18452
rect 16380 18338 16436 18340
rect 16380 18286 16382 18338
rect 16382 18286 16434 18338
rect 16434 18286 16436 18338
rect 16380 18284 16436 18286
rect 16828 18338 16884 18340
rect 16828 18286 16830 18338
rect 16830 18286 16882 18338
rect 16882 18286 16884 18338
rect 16828 18284 16884 18286
rect 16380 17836 16436 17892
rect 16604 17778 16660 17780
rect 16604 17726 16606 17778
rect 16606 17726 16658 17778
rect 16658 17726 16660 17778
rect 16604 17724 16660 17726
rect 17164 17724 17220 17780
rect 17724 20748 17780 20804
rect 17836 20578 17892 20580
rect 17836 20526 17838 20578
rect 17838 20526 17890 20578
rect 17890 20526 17892 20578
rect 17836 20524 17892 20526
rect 18060 20972 18116 21028
rect 17724 20412 17780 20468
rect 17948 20412 18004 20468
rect 17836 20300 17892 20356
rect 17724 20242 17780 20244
rect 17724 20190 17726 20242
rect 17726 20190 17778 20242
rect 17778 20190 17780 20242
rect 17724 20188 17780 20190
rect 18284 21474 18340 21476
rect 18284 21422 18286 21474
rect 18286 21422 18338 21474
rect 18338 21422 18340 21474
rect 18284 21420 18340 21422
rect 18284 21196 18340 21252
rect 17836 19852 17892 19908
rect 17724 19234 17780 19236
rect 17724 19182 17726 19234
rect 17726 19182 17778 19234
rect 17778 19182 17780 19234
rect 17724 19180 17780 19182
rect 17724 18956 17780 19012
rect 17836 18450 17892 18452
rect 17836 18398 17838 18450
rect 17838 18398 17890 18450
rect 17890 18398 17892 18450
rect 17836 18396 17892 18398
rect 18396 20860 18452 20916
rect 18508 21586 18564 21588
rect 18508 21534 18510 21586
rect 18510 21534 18562 21586
rect 18562 21534 18564 21586
rect 18508 21532 18564 21534
rect 18396 20412 18452 20468
rect 18956 22146 19012 22148
rect 18956 22094 18958 22146
rect 18958 22094 19010 22146
rect 19010 22094 19012 22146
rect 18956 22092 19012 22094
rect 18732 21980 18788 22036
rect 18620 21084 18676 21140
rect 18620 20748 18676 20804
rect 18844 20690 18900 20692
rect 18844 20638 18846 20690
rect 18846 20638 18898 20690
rect 18898 20638 18900 20690
rect 18844 20636 18900 20638
rect 18732 19964 18788 20020
rect 19964 26124 20020 26180
rect 22316 26684 22372 26740
rect 23436 31778 23492 31780
rect 23436 31726 23438 31778
rect 23438 31726 23490 31778
rect 23490 31726 23492 31778
rect 23436 31724 23492 31726
rect 23212 31666 23268 31668
rect 23212 31614 23214 31666
rect 23214 31614 23266 31666
rect 23266 31614 23268 31666
rect 23212 31612 23268 31614
rect 23324 31554 23380 31556
rect 23324 31502 23326 31554
rect 23326 31502 23378 31554
rect 23378 31502 23380 31554
rect 23324 31500 23380 31502
rect 24108 32172 24164 32228
rect 24668 31836 24724 31892
rect 24444 31778 24500 31780
rect 24444 31726 24446 31778
rect 24446 31726 24498 31778
rect 24498 31726 24500 31778
rect 24444 31724 24500 31726
rect 23324 30604 23380 30660
rect 25900 37266 25956 37268
rect 25900 37214 25902 37266
rect 25902 37214 25954 37266
rect 25954 37214 25956 37266
rect 25900 37212 25956 37214
rect 25900 36876 25956 36932
rect 26236 36764 26292 36820
rect 25788 35532 25844 35588
rect 26124 36316 26180 36372
rect 26572 36540 26628 36596
rect 26684 35698 26740 35700
rect 26684 35646 26686 35698
rect 26686 35646 26738 35698
rect 26738 35646 26740 35698
rect 26684 35644 26740 35646
rect 28812 38556 28868 38612
rect 28924 38220 28980 38276
rect 30380 38220 30436 38276
rect 27804 37826 27860 37828
rect 27804 37774 27806 37826
rect 27806 37774 27858 37826
rect 27858 37774 27860 37826
rect 27804 37772 27860 37774
rect 27580 37436 27636 37492
rect 28700 37324 28756 37380
rect 27244 36988 27300 37044
rect 27916 37212 27972 37268
rect 27580 36594 27636 36596
rect 27580 36542 27582 36594
rect 27582 36542 27634 36594
rect 27634 36542 27636 36594
rect 27580 36540 27636 36542
rect 27356 35868 27412 35924
rect 25676 34914 25732 34916
rect 25676 34862 25678 34914
rect 25678 34862 25730 34914
rect 25730 34862 25732 34914
rect 25676 34860 25732 34862
rect 26572 34802 26628 34804
rect 26572 34750 26574 34802
rect 26574 34750 26626 34802
rect 26626 34750 26628 34802
rect 26572 34748 26628 34750
rect 25676 34242 25732 34244
rect 25676 34190 25678 34242
rect 25678 34190 25730 34242
rect 25730 34190 25732 34242
rect 25676 34188 25732 34190
rect 26236 34130 26292 34132
rect 26236 34078 26238 34130
rect 26238 34078 26290 34130
rect 26290 34078 26292 34130
rect 26236 34076 26292 34078
rect 26124 34018 26180 34020
rect 26124 33966 26126 34018
rect 26126 33966 26178 34018
rect 26178 33966 26180 34018
rect 26124 33964 26180 33966
rect 26124 33516 26180 33572
rect 26236 33122 26292 33124
rect 26236 33070 26238 33122
rect 26238 33070 26290 33122
rect 26290 33070 26292 33122
rect 26236 33068 26292 33070
rect 26460 33964 26516 34020
rect 26460 33628 26516 33684
rect 25676 31778 25732 31780
rect 25676 31726 25678 31778
rect 25678 31726 25730 31778
rect 25730 31726 25732 31778
rect 25676 31724 25732 31726
rect 26012 31666 26068 31668
rect 26012 31614 26014 31666
rect 26014 31614 26066 31666
rect 26066 31614 26068 31666
rect 26012 31612 26068 31614
rect 22540 29596 22596 29652
rect 22652 27804 22708 27860
rect 22876 27580 22932 27636
rect 22988 27692 23044 27748
rect 20860 26236 20916 26292
rect 19628 25676 19684 25732
rect 19292 25004 19348 25060
rect 19516 24892 19572 24948
rect 20300 25730 20356 25732
rect 20300 25678 20302 25730
rect 20302 25678 20354 25730
rect 20354 25678 20356 25730
rect 20300 25676 20356 25678
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20636 25340 20692 25396
rect 19740 24834 19796 24836
rect 19740 24782 19742 24834
rect 19742 24782 19794 24834
rect 19794 24782 19796 24834
rect 19740 24780 19796 24782
rect 19740 24556 19796 24612
rect 20524 24834 20580 24836
rect 20524 24782 20526 24834
rect 20526 24782 20578 24834
rect 20578 24782 20580 24834
rect 20524 24780 20580 24782
rect 20300 24556 20356 24612
rect 19516 23772 19572 23828
rect 19292 23324 19348 23380
rect 19404 23660 19460 23716
rect 19292 23042 19348 23044
rect 19292 22990 19294 23042
rect 19294 22990 19346 23042
rect 19346 22990 19348 23042
rect 19292 22988 19348 22990
rect 19292 21980 19348 22036
rect 19292 21756 19348 21812
rect 19180 18508 19236 18564
rect 18060 18284 18116 18340
rect 19836 23546 19892 23548
rect 19628 23436 19684 23492
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19628 23212 19684 23268
rect 19964 23324 20020 23380
rect 20412 23212 20468 23268
rect 19964 23042 20020 23044
rect 19964 22990 19966 23042
rect 19966 22990 20018 23042
rect 20018 22990 20020 23042
rect 19964 22988 20020 22990
rect 19964 22092 20020 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19852 21196 19908 21252
rect 20636 23884 20692 23940
rect 20748 23826 20804 23828
rect 20748 23774 20750 23826
rect 20750 23774 20802 23826
rect 20802 23774 20804 23826
rect 20748 23772 20804 23774
rect 20748 23324 20804 23380
rect 22540 26348 22596 26404
rect 21980 25116 22036 25172
rect 21532 24780 21588 24836
rect 20972 23884 21028 23940
rect 21644 24668 21700 24724
rect 21644 23884 21700 23940
rect 21084 23324 21140 23380
rect 20972 23100 21028 23156
rect 20300 21980 20356 22036
rect 21196 22988 21252 23044
rect 22540 25228 22596 25284
rect 22092 24722 22148 24724
rect 22092 24670 22094 24722
rect 22094 24670 22146 24722
rect 22146 24670 22148 24722
rect 22092 24668 22148 24670
rect 22428 25116 22484 25172
rect 21980 23436 22036 23492
rect 22092 23772 22148 23828
rect 21868 23324 21924 23380
rect 21644 23100 21700 23156
rect 21868 23042 21924 23044
rect 21868 22990 21870 23042
rect 21870 22990 21922 23042
rect 21922 22990 21924 23042
rect 21868 22988 21924 22990
rect 21756 22764 21812 22820
rect 19852 20690 19908 20692
rect 19852 20638 19854 20690
rect 19854 20638 19906 20690
rect 19906 20638 19908 20690
rect 19852 20636 19908 20638
rect 20524 22092 20580 22148
rect 20188 20914 20244 20916
rect 20188 20862 20190 20914
rect 20190 20862 20242 20914
rect 20242 20862 20244 20914
rect 20188 20860 20244 20862
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19516 19068 19572 19124
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19404 18172 19460 18228
rect 18956 18060 19012 18116
rect 18396 17778 18452 17780
rect 18396 17726 18398 17778
rect 18398 17726 18450 17778
rect 18450 17726 18452 17778
rect 18396 17724 18452 17726
rect 20748 22146 20804 22148
rect 20748 22094 20750 22146
rect 20750 22094 20802 22146
rect 20802 22094 20804 22146
rect 20748 22092 20804 22094
rect 21868 22540 21924 22596
rect 22428 23938 22484 23940
rect 22428 23886 22430 23938
rect 22430 23886 22482 23938
rect 22482 23886 22484 23938
rect 22428 23884 22484 23886
rect 22204 22540 22260 22596
rect 21420 21756 21476 21812
rect 21532 21980 21588 22036
rect 20748 21644 20804 21700
rect 20524 20860 20580 20916
rect 20860 20636 20916 20692
rect 20412 19292 20468 19348
rect 20300 19010 20356 19012
rect 20300 18958 20302 19010
rect 20302 18958 20354 19010
rect 20354 18958 20356 19010
rect 20300 18956 20356 18958
rect 19740 17836 19796 17892
rect 19292 17724 19348 17780
rect 18172 17612 18228 17668
rect 17052 17276 17108 17332
rect 14812 16994 14868 16996
rect 14812 16942 14814 16994
rect 14814 16942 14866 16994
rect 14866 16942 14868 16994
rect 14812 16940 14868 16942
rect 20412 18172 20468 18228
rect 19852 17724 19908 17780
rect 19964 18060 20020 18116
rect 20412 17890 20468 17892
rect 20412 17838 20414 17890
rect 20414 17838 20466 17890
rect 20466 17838 20468 17890
rect 20412 17836 20468 17838
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 17388 16940 17444 16996
rect 15932 16882 15988 16884
rect 15932 16830 15934 16882
rect 15934 16830 15986 16882
rect 15986 16830 15988 16882
rect 15932 16828 15988 16830
rect 17276 16882 17332 16884
rect 17276 16830 17278 16882
rect 17278 16830 17330 16882
rect 17330 16830 17332 16882
rect 17276 16828 17332 16830
rect 15260 16716 15316 16772
rect 15596 16716 15652 16772
rect 14364 15538 14420 15540
rect 14364 15486 14366 15538
rect 14366 15486 14418 15538
rect 14418 15486 14420 15538
rect 14364 15484 14420 15486
rect 16268 16770 16324 16772
rect 16268 16718 16270 16770
rect 16270 16718 16322 16770
rect 16322 16718 16324 16770
rect 16268 16716 16324 16718
rect 16828 16770 16884 16772
rect 16828 16718 16830 16770
rect 16830 16718 16882 16770
rect 16882 16718 16884 16770
rect 16828 16716 16884 16718
rect 15820 16492 15876 16548
rect 17500 16268 17556 16324
rect 17612 16716 17668 16772
rect 17500 15538 17556 15540
rect 17500 15486 17502 15538
rect 17502 15486 17554 15538
rect 17554 15486 17556 15538
rect 17500 15484 17556 15486
rect 14476 15426 14532 15428
rect 14476 15374 14478 15426
rect 14478 15374 14530 15426
rect 14530 15374 14532 15426
rect 14476 15372 14532 15374
rect 18172 16322 18228 16324
rect 18172 16270 18174 16322
rect 18174 16270 18226 16322
rect 18226 16270 18228 16322
rect 18172 16268 18228 16270
rect 19964 16828 20020 16884
rect 18396 16716 18452 16772
rect 18396 16044 18452 16100
rect 16268 15314 16324 15316
rect 16268 15262 16270 15314
rect 16270 15262 16322 15314
rect 16322 15262 16324 15314
rect 16268 15260 16324 15262
rect 17276 15314 17332 15316
rect 17276 15262 17278 15314
rect 17278 15262 17330 15314
rect 17330 15262 17332 15314
rect 17276 15260 17332 15262
rect 15372 15202 15428 15204
rect 15372 15150 15374 15202
rect 15374 15150 15426 15202
rect 15426 15150 15428 15202
rect 15372 15148 15428 15150
rect 10668 14476 10724 14532
rect 13692 14530 13748 14532
rect 13692 14478 13694 14530
rect 13694 14478 13746 14530
rect 13746 14478 13748 14530
rect 13692 14476 13748 14478
rect 7308 13186 7364 13188
rect 7308 13134 7310 13186
rect 7310 13134 7362 13186
rect 7362 13134 7364 13186
rect 7308 13132 7364 13134
rect 2268 12962 2324 12964
rect 2268 12910 2270 12962
rect 2270 12910 2322 12962
rect 2322 12910 2324 12962
rect 2268 12908 2324 12910
rect 4844 12908 4900 12964
rect 7980 12962 8036 12964
rect 7980 12910 7982 12962
rect 7982 12910 8034 12962
rect 8034 12910 8036 12962
rect 7980 12908 8036 12910
rect 7644 12850 7700 12852
rect 7644 12798 7646 12850
rect 7646 12798 7698 12850
rect 7698 12798 7700 12850
rect 7644 12796 7700 12798
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 5964 11564 6020 11620
rect 6860 11618 6916 11620
rect 6860 11566 6862 11618
rect 6862 11566 6914 11618
rect 6914 11566 6916 11618
rect 6860 11564 6916 11566
rect 8540 12908 8596 12964
rect 8764 12850 8820 12852
rect 8764 12798 8766 12850
rect 8766 12798 8818 12850
rect 8818 12798 8820 12850
rect 8764 12796 8820 12798
rect 8540 12290 8596 12292
rect 8540 12238 8542 12290
rect 8542 12238 8594 12290
rect 8594 12238 8596 12290
rect 8540 12236 8596 12238
rect 16716 15202 16772 15204
rect 16716 15150 16718 15202
rect 16718 15150 16770 15202
rect 16770 15150 16772 15202
rect 16716 15148 16772 15150
rect 18396 15484 18452 15540
rect 18060 15202 18116 15204
rect 18060 15150 18062 15202
rect 18062 15150 18114 15202
rect 18114 15150 18116 15202
rect 18060 15148 18116 15150
rect 19628 16716 19684 16772
rect 18732 16380 18788 16436
rect 19516 16380 19572 16436
rect 18620 16268 18676 16324
rect 19404 16210 19460 16212
rect 19404 16158 19406 16210
rect 19406 16158 19458 16210
rect 19458 16158 19460 16210
rect 19404 16156 19460 16158
rect 19292 16098 19348 16100
rect 19292 16046 19294 16098
rect 19294 16046 19346 16098
rect 19346 16046 19348 16098
rect 19292 16044 19348 16046
rect 19180 15372 19236 15428
rect 18732 15148 18788 15204
rect 14252 14476 14308 14532
rect 14924 14530 14980 14532
rect 14924 14478 14926 14530
rect 14926 14478 14978 14530
rect 14978 14478 14980 14530
rect 14924 14476 14980 14478
rect 10892 13074 10948 13076
rect 10892 13022 10894 13074
rect 10894 13022 10946 13074
rect 10946 13022 10948 13074
rect 10892 13020 10948 13022
rect 12012 13074 12068 13076
rect 12012 13022 12014 13074
rect 12014 13022 12066 13074
rect 12066 13022 12068 13074
rect 12012 13020 12068 13022
rect 9996 12236 10052 12292
rect 11228 12684 11284 12740
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 9660 11170 9716 11172
rect 9660 11118 9662 11170
rect 9662 11118 9714 11170
rect 9714 11118 9716 11170
rect 9660 11116 9716 11118
rect 10780 11282 10836 11284
rect 10780 11230 10782 11282
rect 10782 11230 10834 11282
rect 10834 11230 10836 11282
rect 10780 11228 10836 11230
rect 10332 11116 10388 11172
rect 9436 9996 9492 10052
rect 10780 10050 10836 10052
rect 10780 9998 10782 10050
rect 10782 9998 10834 10050
rect 10834 9998 10836 10050
rect 10780 9996 10836 9998
rect 11340 11900 11396 11956
rect 11900 12738 11956 12740
rect 11900 12686 11902 12738
rect 11902 12686 11954 12738
rect 11954 12686 11956 12738
rect 11900 12684 11956 12686
rect 14700 13020 14756 13076
rect 13580 11900 13636 11956
rect 12908 11506 12964 11508
rect 12908 11454 12910 11506
rect 12910 11454 12962 11506
rect 12962 11454 12964 11506
rect 12908 11452 12964 11454
rect 14364 11452 14420 11508
rect 11452 10444 11508 10500
rect 12460 10498 12516 10500
rect 12460 10446 12462 10498
rect 12462 10446 12514 10498
rect 12514 10446 12516 10498
rect 12460 10444 12516 10446
rect 12572 9938 12628 9940
rect 12572 9886 12574 9938
rect 12574 9886 12626 9938
rect 12626 9886 12628 9938
rect 12572 9884 12628 9886
rect 13020 9938 13076 9940
rect 13020 9886 13022 9938
rect 13022 9886 13074 9938
rect 13074 9886 13076 9938
rect 13020 9884 13076 9886
rect 13692 9938 13748 9940
rect 13692 9886 13694 9938
rect 13694 9886 13746 9938
rect 13746 9886 13748 9938
rect 13692 9884 13748 9886
rect 13916 11228 13972 11284
rect 15932 13916 15988 13972
rect 16828 13970 16884 13972
rect 16828 13918 16830 13970
rect 16830 13918 16882 13970
rect 16882 13918 16884 13970
rect 16828 13916 16884 13918
rect 16380 13858 16436 13860
rect 16380 13806 16382 13858
rect 16382 13806 16434 13858
rect 16434 13806 16436 13858
rect 16380 13804 16436 13806
rect 20188 16044 20244 16100
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19628 15314 19684 15316
rect 19628 15262 19630 15314
rect 19630 15262 19682 15314
rect 19682 15262 19684 15314
rect 19628 15260 19684 15262
rect 19740 15148 19796 15204
rect 18508 14924 18564 14980
rect 17836 13858 17892 13860
rect 17836 13806 17838 13858
rect 17838 13806 17890 13858
rect 17890 13806 17892 13858
rect 17836 13804 17892 13806
rect 19068 15036 19124 15092
rect 19068 14812 19124 14868
rect 19292 14588 19348 14644
rect 18844 13468 18900 13524
rect 15260 13074 15316 13076
rect 15260 13022 15262 13074
rect 15262 13022 15314 13074
rect 15314 13022 15316 13074
rect 15260 13020 15316 13022
rect 15596 13020 15652 13076
rect 18508 13074 18564 13076
rect 18508 13022 18510 13074
rect 18510 13022 18562 13074
rect 18562 13022 18564 13074
rect 18508 13020 18564 13022
rect 18508 12850 18564 12852
rect 18508 12798 18510 12850
rect 18510 12798 18562 12850
rect 18562 12798 18564 12850
rect 18508 12796 18564 12798
rect 19292 13468 19348 13524
rect 21420 19122 21476 19124
rect 21420 19070 21422 19122
rect 21422 19070 21474 19122
rect 21474 19070 21476 19122
rect 21420 19068 21476 19070
rect 21308 19010 21364 19012
rect 21308 18958 21310 19010
rect 21310 18958 21362 19010
rect 21362 18958 21364 19010
rect 21308 18956 21364 18958
rect 21420 18338 21476 18340
rect 21420 18286 21422 18338
rect 21422 18286 21474 18338
rect 21474 18286 21476 18338
rect 21420 18284 21476 18286
rect 21196 17948 21252 18004
rect 20748 17724 20804 17780
rect 20748 17388 20804 17444
rect 21084 16156 21140 16212
rect 20524 16044 20580 16100
rect 20860 15260 20916 15316
rect 21308 17836 21364 17892
rect 22204 22146 22260 22148
rect 22204 22094 22206 22146
rect 22206 22094 22258 22146
rect 22258 22094 22260 22146
rect 22204 22092 22260 22094
rect 22428 21644 22484 21700
rect 22204 20972 22260 21028
rect 22988 26684 23044 26740
rect 22652 25004 22708 25060
rect 23212 26402 23268 26404
rect 23212 26350 23214 26402
rect 23214 26350 23266 26402
rect 23266 26350 23268 26402
rect 23212 26348 23268 26350
rect 22988 25676 23044 25732
rect 22876 25506 22932 25508
rect 22876 25454 22878 25506
rect 22878 25454 22930 25506
rect 22930 25454 22932 25506
rect 22876 25452 22932 25454
rect 26124 31218 26180 31220
rect 26124 31166 26126 31218
rect 26126 31166 26178 31218
rect 26178 31166 26180 31218
rect 26124 31164 26180 31166
rect 26012 30994 26068 30996
rect 26012 30942 26014 30994
rect 26014 30942 26066 30994
rect 26066 30942 26068 30994
rect 26012 30940 26068 30942
rect 25900 30156 25956 30212
rect 24220 29932 24276 29988
rect 24220 29708 24276 29764
rect 24556 30044 24612 30100
rect 25004 30098 25060 30100
rect 25004 30046 25006 30098
rect 25006 30046 25058 30098
rect 25058 30046 25060 30098
rect 25004 30044 25060 30046
rect 24668 29932 24724 29988
rect 23772 28082 23828 28084
rect 23772 28030 23774 28082
rect 23774 28030 23826 28082
rect 23826 28030 23828 28082
rect 23772 28028 23828 28030
rect 23436 26290 23492 26292
rect 23436 26238 23438 26290
rect 23438 26238 23490 26290
rect 23490 26238 23492 26290
rect 23436 26236 23492 26238
rect 22988 24834 23044 24836
rect 22988 24782 22990 24834
rect 22990 24782 23042 24834
rect 23042 24782 23044 24834
rect 22988 24780 23044 24782
rect 22652 23772 22708 23828
rect 21756 20690 21812 20692
rect 21756 20638 21758 20690
rect 21758 20638 21810 20690
rect 21810 20638 21812 20690
rect 21756 20636 21812 20638
rect 22092 20524 22148 20580
rect 22204 19346 22260 19348
rect 22204 19294 22206 19346
rect 22206 19294 22258 19346
rect 22258 19294 22260 19346
rect 22204 19292 22260 19294
rect 21644 18450 21700 18452
rect 21644 18398 21646 18450
rect 21646 18398 21698 18450
rect 21698 18398 21700 18450
rect 21644 18396 21700 18398
rect 21532 17500 21588 17556
rect 21532 17276 21588 17332
rect 21644 18060 21700 18116
rect 21308 16098 21364 16100
rect 21308 16046 21310 16098
rect 21310 16046 21362 16098
rect 21362 16046 21364 16098
rect 21308 16044 21364 16046
rect 21196 15820 21252 15876
rect 21980 18338 22036 18340
rect 21980 18286 21982 18338
rect 21982 18286 22034 18338
rect 22034 18286 22036 18338
rect 21980 18284 22036 18286
rect 21868 17612 21924 17668
rect 21980 16882 22036 16884
rect 21980 16830 21982 16882
rect 21982 16830 22034 16882
rect 22034 16830 22036 16882
rect 21980 16828 22036 16830
rect 22652 20802 22708 20804
rect 22652 20750 22654 20802
rect 22654 20750 22706 20802
rect 22706 20750 22708 20802
rect 22652 20748 22708 20750
rect 22876 23324 22932 23380
rect 22876 22764 22932 22820
rect 23884 26236 23940 26292
rect 23772 26178 23828 26180
rect 23772 26126 23774 26178
rect 23774 26126 23826 26178
rect 23826 26126 23828 26178
rect 23772 26124 23828 26126
rect 23996 26124 24052 26180
rect 23772 25618 23828 25620
rect 23772 25566 23774 25618
rect 23774 25566 23826 25618
rect 23826 25566 23828 25618
rect 23772 25564 23828 25566
rect 24220 25676 24276 25732
rect 23660 25452 23716 25508
rect 23324 25116 23380 25172
rect 25788 29986 25844 29988
rect 25788 29934 25790 29986
rect 25790 29934 25842 29986
rect 25842 29934 25844 29986
rect 25788 29932 25844 29934
rect 25564 29372 25620 29428
rect 25116 28028 25172 28084
rect 24780 27804 24836 27860
rect 24780 27132 24836 27188
rect 25228 29314 25284 29316
rect 25228 29262 25230 29314
rect 25230 29262 25282 29314
rect 25282 29262 25284 29314
rect 25228 29260 25284 29262
rect 25340 29202 25396 29204
rect 25340 29150 25342 29202
rect 25342 29150 25394 29202
rect 25394 29150 25396 29202
rect 25340 29148 25396 29150
rect 25340 27746 25396 27748
rect 25340 27694 25342 27746
rect 25342 27694 25394 27746
rect 25394 27694 25396 27746
rect 25340 27692 25396 27694
rect 25452 27186 25508 27188
rect 25452 27134 25454 27186
rect 25454 27134 25506 27186
rect 25506 27134 25508 27186
rect 25452 27132 25508 27134
rect 25228 25506 25284 25508
rect 25228 25454 25230 25506
rect 25230 25454 25282 25506
rect 25282 25454 25284 25506
rect 25228 25452 25284 25454
rect 24444 25340 24500 25396
rect 24444 25116 24500 25172
rect 23996 24722 24052 24724
rect 23996 24670 23998 24722
rect 23998 24670 24050 24722
rect 24050 24670 24052 24722
rect 23996 24668 24052 24670
rect 23772 24556 23828 24612
rect 23212 23884 23268 23940
rect 23996 23938 24052 23940
rect 23996 23886 23998 23938
rect 23998 23886 24050 23938
rect 24050 23886 24052 23938
rect 23996 23884 24052 23886
rect 25228 24668 25284 24724
rect 25004 24556 25060 24612
rect 24332 23772 24388 23828
rect 22876 20914 22932 20916
rect 22876 20862 22878 20914
rect 22878 20862 22930 20914
rect 22930 20862 22932 20914
rect 22876 20860 22932 20862
rect 23100 22482 23156 22484
rect 23100 22430 23102 22482
rect 23102 22430 23154 22482
rect 23154 22430 23156 22482
rect 23100 22428 23156 22430
rect 24220 22988 24276 23044
rect 24556 23154 24612 23156
rect 24556 23102 24558 23154
rect 24558 23102 24610 23154
rect 24610 23102 24612 23154
rect 24556 23100 24612 23102
rect 24444 22316 24500 22372
rect 23660 21644 23716 21700
rect 23548 21196 23604 21252
rect 23324 20972 23380 21028
rect 23660 20578 23716 20580
rect 23660 20526 23662 20578
rect 23662 20526 23714 20578
rect 23714 20526 23716 20578
rect 23660 20524 23716 20526
rect 23772 20636 23828 20692
rect 22988 20300 23044 20356
rect 22764 19852 22820 19908
rect 22428 17948 22484 18004
rect 22764 17666 22820 17668
rect 22764 17614 22766 17666
rect 22766 17614 22818 17666
rect 22818 17614 22820 17666
rect 22764 17612 22820 17614
rect 22988 18284 23044 18340
rect 23212 17948 23268 18004
rect 22988 17052 23044 17108
rect 22428 16828 22484 16884
rect 20188 14530 20244 14532
rect 20188 14478 20190 14530
rect 20190 14478 20242 14530
rect 20242 14478 20244 14530
rect 20188 14476 20244 14478
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20412 13074 20468 13076
rect 20412 13022 20414 13074
rect 20414 13022 20466 13074
rect 20466 13022 20468 13074
rect 20412 13020 20468 13022
rect 20524 12908 20580 12964
rect 16716 11676 16772 11732
rect 15372 9938 15428 9940
rect 15372 9886 15374 9938
rect 15374 9886 15426 9938
rect 15426 9886 15428 9938
rect 15372 9884 15428 9886
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 18060 11452 18116 11508
rect 18732 11452 18788 11508
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 18172 3612 18228 3668
rect 18844 9884 18900 9940
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 20300 12236 20356 12292
rect 19964 11900 20020 11956
rect 19852 11788 19908 11844
rect 20412 11788 20468 11844
rect 19628 11676 19684 11732
rect 21308 14924 21364 14980
rect 21532 14700 21588 14756
rect 21644 14418 21700 14420
rect 21644 14366 21646 14418
rect 21646 14366 21698 14418
rect 21698 14366 21700 14418
rect 21644 14364 21700 14366
rect 21308 13804 21364 13860
rect 21420 13634 21476 13636
rect 21420 13582 21422 13634
rect 21422 13582 21474 13634
rect 21474 13582 21476 13634
rect 21420 13580 21476 13582
rect 21868 14700 21924 14756
rect 22092 15314 22148 15316
rect 22092 15262 22094 15314
rect 22094 15262 22146 15314
rect 22146 15262 22148 15314
rect 22092 15260 22148 15262
rect 22204 14530 22260 14532
rect 22204 14478 22206 14530
rect 22206 14478 22258 14530
rect 22258 14478 22260 14530
rect 22204 14476 22260 14478
rect 23100 17276 23156 17332
rect 23324 15314 23380 15316
rect 23324 15262 23326 15314
rect 23326 15262 23378 15314
rect 23378 15262 23380 15314
rect 23324 15260 23380 15262
rect 22540 14588 22596 14644
rect 21084 12908 21140 12964
rect 21868 12796 21924 12852
rect 20860 12178 20916 12180
rect 20860 12126 20862 12178
rect 20862 12126 20914 12178
rect 20914 12126 20916 12178
rect 20860 12124 20916 12126
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19740 10050 19796 10052
rect 19740 9998 19742 10050
rect 19742 9998 19794 10050
rect 19794 9998 19796 10050
rect 19740 9996 19796 9998
rect 20972 11228 21028 11284
rect 20972 9996 21028 10052
rect 20748 9826 20804 9828
rect 20748 9774 20750 9826
rect 20750 9774 20802 9826
rect 20802 9774 20804 9826
rect 20748 9772 20804 9774
rect 19628 9548 19684 9604
rect 20524 9714 20580 9716
rect 20524 9662 20526 9714
rect 20526 9662 20578 9714
rect 20578 9662 20580 9714
rect 20524 9660 20580 9662
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 18844 3666 18900 3668
rect 18844 3614 18846 3666
rect 18846 3614 18898 3666
rect 18898 3614 18900 3666
rect 18844 3612 18900 3614
rect 22092 12962 22148 12964
rect 22092 12910 22094 12962
rect 22094 12910 22146 12962
rect 22146 12910 22148 12962
rect 22092 12908 22148 12910
rect 21868 11282 21924 11284
rect 21868 11230 21870 11282
rect 21870 11230 21922 11282
rect 21922 11230 21924 11282
rect 21868 11228 21924 11230
rect 22428 13916 22484 13972
rect 22652 12796 22708 12852
rect 22204 12178 22260 12180
rect 22204 12126 22206 12178
rect 22206 12126 22258 12178
rect 22258 12126 22260 12178
rect 22204 12124 22260 12126
rect 22204 10498 22260 10500
rect 22204 10446 22206 10498
rect 22206 10446 22258 10498
rect 22258 10446 22260 10498
rect 22204 10444 22260 10446
rect 21644 9938 21700 9940
rect 21644 9886 21646 9938
rect 21646 9886 21698 9938
rect 21698 9886 21700 9938
rect 21644 9884 21700 9886
rect 21308 9826 21364 9828
rect 21308 9774 21310 9826
rect 21310 9774 21362 9826
rect 21362 9774 21364 9826
rect 21308 9772 21364 9774
rect 21868 9772 21924 9828
rect 21420 9548 21476 9604
rect 24220 21362 24276 21364
rect 24220 21310 24222 21362
rect 24222 21310 24274 21362
rect 24274 21310 24276 21362
rect 24220 21308 24276 21310
rect 24220 20914 24276 20916
rect 24220 20862 24222 20914
rect 24222 20862 24274 20914
rect 24274 20862 24276 20914
rect 24220 20860 24276 20862
rect 23996 20802 24052 20804
rect 23996 20750 23998 20802
rect 23998 20750 24050 20802
rect 24050 20750 24052 20802
rect 23996 20748 24052 20750
rect 23996 20188 24052 20244
rect 24108 19628 24164 19684
rect 24220 20300 24276 20356
rect 24108 19234 24164 19236
rect 24108 19182 24110 19234
rect 24110 19182 24162 19234
rect 24162 19182 24164 19234
rect 24108 19180 24164 19182
rect 24668 21084 24724 21140
rect 24780 22988 24836 23044
rect 25452 25340 25508 25396
rect 26012 29708 26068 29764
rect 25788 29314 25844 29316
rect 25788 29262 25790 29314
rect 25790 29262 25842 29314
rect 25842 29262 25844 29314
rect 25788 29260 25844 29262
rect 25900 29148 25956 29204
rect 25900 27074 25956 27076
rect 25900 27022 25902 27074
rect 25902 27022 25954 27074
rect 25954 27022 25956 27074
rect 25900 27020 25956 27022
rect 25564 25228 25620 25284
rect 25900 24946 25956 24948
rect 25900 24894 25902 24946
rect 25902 24894 25954 24946
rect 25954 24894 25956 24946
rect 25900 24892 25956 24894
rect 25900 24668 25956 24724
rect 26348 31890 26404 31892
rect 26348 31838 26350 31890
rect 26350 31838 26402 31890
rect 26402 31838 26404 31890
rect 26348 31836 26404 31838
rect 26572 31778 26628 31780
rect 26572 31726 26574 31778
rect 26574 31726 26626 31778
rect 26626 31726 26628 31778
rect 26572 31724 26628 31726
rect 27692 36370 27748 36372
rect 27692 36318 27694 36370
rect 27694 36318 27746 36370
rect 27746 36318 27748 36370
rect 27692 36316 27748 36318
rect 28476 36370 28532 36372
rect 28476 36318 28478 36370
rect 28478 36318 28530 36370
rect 28530 36318 28532 36370
rect 28476 36316 28532 36318
rect 26908 34636 26964 34692
rect 27356 34690 27412 34692
rect 27356 34638 27358 34690
rect 27358 34638 27410 34690
rect 27410 34638 27412 34690
rect 27356 34636 27412 34638
rect 27244 34300 27300 34356
rect 27132 34130 27188 34132
rect 27132 34078 27134 34130
rect 27134 34078 27186 34130
rect 27186 34078 27188 34130
rect 27132 34076 27188 34078
rect 27132 33852 27188 33908
rect 27356 33740 27412 33796
rect 26908 32674 26964 32676
rect 26908 32622 26910 32674
rect 26910 32622 26962 32674
rect 26962 32622 26964 32674
rect 26908 32620 26964 32622
rect 27020 31836 27076 31892
rect 26796 31724 26852 31780
rect 26908 31666 26964 31668
rect 26908 31614 26910 31666
rect 26910 31614 26962 31666
rect 26962 31614 26964 31666
rect 26908 31612 26964 31614
rect 26796 31164 26852 31220
rect 26684 30940 26740 30996
rect 26348 30098 26404 30100
rect 26348 30046 26350 30098
rect 26350 30046 26402 30098
rect 26402 30046 26404 30098
rect 26348 30044 26404 30046
rect 26572 30044 26628 30100
rect 26348 29426 26404 29428
rect 26348 29374 26350 29426
rect 26350 29374 26402 29426
rect 26402 29374 26404 29426
rect 26348 29372 26404 29374
rect 26348 28252 26404 28308
rect 26236 27074 26292 27076
rect 26236 27022 26238 27074
rect 26238 27022 26290 27074
rect 26290 27022 26292 27074
rect 26236 27020 26292 27022
rect 27356 33068 27412 33124
rect 27356 32396 27412 32452
rect 28364 35922 28420 35924
rect 28364 35870 28366 35922
rect 28366 35870 28418 35922
rect 28418 35870 28420 35922
rect 28364 35868 28420 35870
rect 27916 35586 27972 35588
rect 27916 35534 27918 35586
rect 27918 35534 27970 35586
rect 27970 35534 27972 35586
rect 27916 35532 27972 35534
rect 27916 34300 27972 34356
rect 28364 34636 28420 34692
rect 28028 34188 28084 34244
rect 28140 34076 28196 34132
rect 27804 33516 27860 33572
rect 27916 33740 27972 33796
rect 27692 31836 27748 31892
rect 28028 32674 28084 32676
rect 28028 32622 28030 32674
rect 28030 32622 28082 32674
rect 28082 32622 28084 32674
rect 28028 32620 28084 32622
rect 28140 32396 28196 32452
rect 27804 31724 27860 31780
rect 28028 31890 28084 31892
rect 28028 31838 28030 31890
rect 28030 31838 28082 31890
rect 28082 31838 28084 31890
rect 28028 31836 28084 31838
rect 28252 31724 28308 31780
rect 27580 31666 27636 31668
rect 27580 31614 27582 31666
rect 27582 31614 27634 31666
rect 27634 31614 27636 31666
rect 27580 31612 27636 31614
rect 27244 31500 27300 31556
rect 27468 30882 27524 30884
rect 27468 30830 27470 30882
rect 27470 30830 27522 30882
rect 27522 30830 27524 30882
rect 27468 30828 27524 30830
rect 27916 30210 27972 30212
rect 27916 30158 27918 30210
rect 27918 30158 27970 30210
rect 27970 30158 27972 30210
rect 27916 30156 27972 30158
rect 26908 30098 26964 30100
rect 26908 30046 26910 30098
rect 26910 30046 26962 30098
rect 26962 30046 26964 30098
rect 26908 30044 26964 30046
rect 27804 30044 27860 30100
rect 27356 28754 27412 28756
rect 27356 28702 27358 28754
rect 27358 28702 27410 28754
rect 27410 28702 27412 28754
rect 27356 28700 27412 28702
rect 26572 27858 26628 27860
rect 26572 27806 26574 27858
rect 26574 27806 26626 27858
rect 26626 27806 26628 27858
rect 26572 27804 26628 27806
rect 26684 27692 26740 27748
rect 27020 28530 27076 28532
rect 27020 28478 27022 28530
rect 27022 28478 27074 28530
rect 27074 28478 27076 28530
rect 27020 28476 27076 28478
rect 27804 28530 27860 28532
rect 27804 28478 27806 28530
rect 27806 28478 27858 28530
rect 27858 28478 27860 28530
rect 27804 28476 27860 28478
rect 27580 27804 27636 27860
rect 26684 27356 26740 27412
rect 27468 27186 27524 27188
rect 27468 27134 27470 27186
rect 27470 27134 27522 27186
rect 27522 27134 27524 27186
rect 27468 27132 27524 27134
rect 26460 26796 26516 26852
rect 26236 26460 26292 26516
rect 26684 26124 26740 26180
rect 27356 26236 27412 26292
rect 26012 23772 26068 23828
rect 25676 22988 25732 23044
rect 26236 23042 26292 23044
rect 26236 22990 26238 23042
rect 26238 22990 26290 23042
rect 26290 22990 26292 23042
rect 26236 22988 26292 22990
rect 25900 22930 25956 22932
rect 25900 22878 25902 22930
rect 25902 22878 25954 22930
rect 25954 22878 25956 22930
rect 25900 22876 25956 22878
rect 25788 22370 25844 22372
rect 25788 22318 25790 22370
rect 25790 22318 25842 22370
rect 25842 22318 25844 22370
rect 25788 22316 25844 22318
rect 25452 22092 25508 22148
rect 24444 20524 24500 20580
rect 25340 21810 25396 21812
rect 25340 21758 25342 21810
rect 25342 21758 25394 21810
rect 25394 21758 25396 21810
rect 25340 21756 25396 21758
rect 25452 21196 25508 21252
rect 25228 20242 25284 20244
rect 25228 20190 25230 20242
rect 25230 20190 25282 20242
rect 25282 20190 25284 20242
rect 25228 20188 25284 20190
rect 24780 20018 24836 20020
rect 24780 19966 24782 20018
rect 24782 19966 24834 20018
rect 24834 19966 24836 20018
rect 24780 19964 24836 19966
rect 24556 19794 24612 19796
rect 24556 19742 24558 19794
rect 24558 19742 24610 19794
rect 24610 19742 24612 19794
rect 24556 19740 24612 19742
rect 25452 20076 25508 20132
rect 24332 19404 24388 19460
rect 24668 19516 24724 19572
rect 23660 17948 23716 18004
rect 23772 18172 23828 18228
rect 25340 19458 25396 19460
rect 25340 19406 25342 19458
rect 25342 19406 25394 19458
rect 25394 19406 25396 19458
rect 25340 19404 25396 19406
rect 24892 19122 24948 19124
rect 24892 19070 24894 19122
rect 24894 19070 24946 19122
rect 24946 19070 24948 19122
rect 24892 19068 24948 19070
rect 24556 18060 24612 18116
rect 24108 17948 24164 18004
rect 24556 16994 24612 16996
rect 24556 16942 24558 16994
rect 24558 16942 24610 16994
rect 24610 16942 24612 16994
rect 24556 16940 24612 16942
rect 23996 16044 24052 16100
rect 26012 21084 26068 21140
rect 25788 20412 25844 20468
rect 25676 19234 25732 19236
rect 25676 19182 25678 19234
rect 25678 19182 25730 19234
rect 25730 19182 25732 19234
rect 25676 19180 25732 19182
rect 25900 19180 25956 19236
rect 26236 20130 26292 20132
rect 26236 20078 26238 20130
rect 26238 20078 26290 20130
rect 26290 20078 26292 20130
rect 26236 20076 26292 20078
rect 26236 19852 26292 19908
rect 26124 19404 26180 19460
rect 26796 25452 26852 25508
rect 27244 24834 27300 24836
rect 27244 24782 27246 24834
rect 27246 24782 27298 24834
rect 27298 24782 27300 24834
rect 27244 24780 27300 24782
rect 26684 24668 26740 24724
rect 28140 26962 28196 26964
rect 28140 26910 28142 26962
rect 28142 26910 28194 26962
rect 28194 26910 28196 26962
rect 28140 26908 28196 26910
rect 29484 37324 29540 37380
rect 30268 37436 30324 37492
rect 29036 36876 29092 36932
rect 29820 37266 29876 37268
rect 29820 37214 29822 37266
rect 29822 37214 29874 37266
rect 29874 37214 29876 37266
rect 29820 37212 29876 37214
rect 29820 36876 29876 36932
rect 29708 36482 29764 36484
rect 29708 36430 29710 36482
rect 29710 36430 29762 36482
rect 29762 36430 29764 36482
rect 29708 36428 29764 36430
rect 29596 36316 29652 36372
rect 29372 36204 29428 36260
rect 30268 36204 30324 36260
rect 28812 35586 28868 35588
rect 28812 35534 28814 35586
rect 28814 35534 28866 35586
rect 28866 35534 28868 35586
rect 28812 35532 28868 35534
rect 30268 35586 30324 35588
rect 30268 35534 30270 35586
rect 30270 35534 30322 35586
rect 30322 35534 30324 35586
rect 30268 35532 30324 35534
rect 28476 32620 28532 32676
rect 28588 31666 28644 31668
rect 28588 31614 28590 31666
rect 28590 31614 28642 31666
rect 28642 31614 28644 31666
rect 28588 31612 28644 31614
rect 28588 29484 28644 29540
rect 28588 27804 28644 27860
rect 30716 36428 30772 36484
rect 30940 36316 30996 36372
rect 30828 36204 30884 36260
rect 30492 35532 30548 35588
rect 29820 34860 29876 34916
rect 29372 34690 29428 34692
rect 29372 34638 29374 34690
rect 29374 34638 29426 34690
rect 29426 34638 29428 34690
rect 29372 34636 29428 34638
rect 29372 34354 29428 34356
rect 29372 34302 29374 34354
rect 29374 34302 29426 34354
rect 29426 34302 29428 34354
rect 29372 34300 29428 34302
rect 30828 35644 30884 35700
rect 31612 37436 31668 37492
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 31836 37436 31892 37492
rect 32396 37490 32452 37492
rect 32396 37438 32398 37490
rect 32398 37438 32450 37490
rect 32450 37438 32452 37490
rect 32396 37436 32452 37438
rect 31388 37378 31444 37380
rect 31388 37326 31390 37378
rect 31390 37326 31442 37378
rect 31442 37326 31444 37378
rect 31388 37324 31444 37326
rect 32732 37324 32788 37380
rect 31500 37266 31556 37268
rect 31500 37214 31502 37266
rect 31502 37214 31554 37266
rect 31554 37214 31556 37266
rect 31500 37212 31556 37214
rect 31276 36876 31332 36932
rect 34972 37490 35028 37492
rect 34972 37438 34974 37490
rect 34974 37438 35026 37490
rect 35026 37438 35028 37490
rect 34972 37436 35028 37438
rect 33740 37324 33796 37380
rect 33628 37266 33684 37268
rect 33628 37214 33630 37266
rect 33630 37214 33682 37266
rect 33682 37214 33684 37266
rect 33628 37212 33684 37214
rect 32508 36876 32564 36932
rect 32060 36428 32116 36484
rect 31948 36370 32004 36372
rect 31948 36318 31950 36370
rect 31950 36318 32002 36370
rect 32002 36318 32004 36370
rect 31948 36316 32004 36318
rect 32060 35698 32116 35700
rect 32060 35646 32062 35698
rect 32062 35646 32114 35698
rect 32114 35646 32116 35698
rect 32060 35644 32116 35646
rect 30828 34860 30884 34916
rect 31388 34914 31444 34916
rect 31388 34862 31390 34914
rect 31390 34862 31442 34914
rect 31442 34862 31444 34914
rect 31388 34860 31444 34862
rect 30940 34690 30996 34692
rect 30940 34638 30942 34690
rect 30942 34638 30994 34690
rect 30994 34638 30996 34690
rect 30940 34636 30996 34638
rect 30828 34354 30884 34356
rect 30828 34302 30830 34354
rect 30830 34302 30882 34354
rect 30882 34302 30884 34354
rect 30828 34300 30884 34302
rect 29820 34076 29876 34132
rect 30492 34130 30548 34132
rect 30492 34078 30494 34130
rect 30494 34078 30546 34130
rect 30546 34078 30548 34130
rect 30492 34076 30548 34078
rect 29148 31778 29204 31780
rect 29148 31726 29150 31778
rect 29150 31726 29202 31778
rect 29202 31726 29204 31778
rect 29148 31724 29204 31726
rect 29260 31666 29316 31668
rect 29260 31614 29262 31666
rect 29262 31614 29314 31666
rect 29314 31614 29316 31666
rect 29260 31612 29316 31614
rect 29260 30828 29316 30884
rect 29148 30210 29204 30212
rect 29148 30158 29150 30210
rect 29150 30158 29202 30210
rect 29202 30158 29204 30210
rect 29148 30156 29204 30158
rect 30380 33628 30436 33684
rect 30492 33234 30548 33236
rect 30492 33182 30494 33234
rect 30494 33182 30546 33234
rect 30546 33182 30548 33234
rect 30492 33180 30548 33182
rect 30828 32786 30884 32788
rect 30828 32734 30830 32786
rect 30830 32734 30882 32786
rect 30882 32734 30884 32786
rect 30828 32732 30884 32734
rect 30492 31836 30548 31892
rect 29820 31666 29876 31668
rect 29820 31614 29822 31666
rect 29822 31614 29874 31666
rect 29874 31614 29876 31666
rect 29820 31612 29876 31614
rect 30604 31666 30660 31668
rect 30604 31614 30606 31666
rect 30606 31614 30658 31666
rect 30658 31614 30660 31666
rect 30604 31612 30660 31614
rect 31836 34690 31892 34692
rect 31836 34638 31838 34690
rect 31838 34638 31890 34690
rect 31890 34638 31892 34690
rect 31836 34636 31892 34638
rect 31500 33346 31556 33348
rect 31500 33294 31502 33346
rect 31502 33294 31554 33346
rect 31554 33294 31556 33346
rect 31500 33292 31556 33294
rect 30940 32060 30996 32116
rect 30940 31890 30996 31892
rect 30940 31838 30942 31890
rect 30942 31838 30994 31890
rect 30994 31838 30996 31890
rect 30940 31836 30996 31838
rect 31500 32060 31556 32116
rect 31388 31836 31444 31892
rect 30716 31388 30772 31444
rect 32844 36876 32900 36932
rect 32060 33852 32116 33908
rect 32172 33292 32228 33348
rect 32396 33628 32452 33684
rect 32508 33852 32564 33908
rect 32508 33404 32564 33460
rect 32284 33234 32340 33236
rect 32284 33182 32286 33234
rect 32286 33182 32338 33234
rect 32338 33182 32340 33234
rect 32284 33180 32340 33182
rect 31724 31948 31780 32004
rect 32508 31948 32564 32004
rect 32060 31836 32116 31892
rect 31836 31778 31892 31780
rect 31836 31726 31838 31778
rect 31838 31726 31890 31778
rect 31890 31726 31892 31778
rect 31836 31724 31892 31726
rect 31612 31612 31668 31668
rect 31164 31388 31220 31444
rect 31500 31388 31556 31444
rect 31612 31218 31668 31220
rect 31612 31166 31614 31218
rect 31614 31166 31666 31218
rect 31666 31166 31668 31218
rect 31612 31164 31668 31166
rect 32172 31052 32228 31108
rect 30604 30716 30660 30772
rect 29596 29820 29652 29876
rect 28700 27356 28756 27412
rect 29148 28642 29204 28644
rect 29148 28590 29150 28642
rect 29150 28590 29202 28642
rect 29202 28590 29204 28642
rect 29148 28588 29204 28590
rect 28364 26236 28420 26292
rect 29036 26796 29092 26852
rect 27692 26124 27748 26180
rect 26684 23772 26740 23828
rect 26460 23154 26516 23156
rect 26460 23102 26462 23154
rect 26462 23102 26514 23154
rect 26514 23102 26516 23154
rect 26460 23100 26516 23102
rect 26796 22988 26852 23044
rect 28140 24892 28196 24948
rect 28252 25004 28308 25060
rect 30380 29260 30436 29316
rect 29820 28588 29876 28644
rect 30380 28642 30436 28644
rect 30380 28590 30382 28642
rect 30382 28590 30434 28642
rect 30434 28590 30436 28642
rect 30380 28588 30436 28590
rect 29708 28082 29764 28084
rect 29708 28030 29710 28082
rect 29710 28030 29762 28082
rect 29762 28030 29764 28082
rect 29708 28028 29764 28030
rect 29596 27804 29652 27860
rect 30380 27858 30436 27860
rect 30380 27806 30382 27858
rect 30382 27806 30434 27858
rect 30434 27806 30436 27858
rect 30380 27804 30436 27806
rect 30716 28700 30772 28756
rect 30828 29596 30884 29652
rect 30716 28082 30772 28084
rect 30716 28030 30718 28082
rect 30718 28030 30770 28082
rect 30770 28030 30772 28082
rect 30716 28028 30772 28030
rect 30940 28028 30996 28084
rect 31052 28476 31108 28532
rect 30604 27692 30660 27748
rect 29820 27132 29876 27188
rect 29484 27020 29540 27076
rect 29260 26962 29316 26964
rect 29260 26910 29262 26962
rect 29262 26910 29314 26962
rect 29314 26910 29316 26962
rect 29260 26908 29316 26910
rect 29148 26124 29204 26180
rect 28812 25452 28868 25508
rect 28476 24780 28532 24836
rect 29484 26124 29540 26180
rect 30940 26796 30996 26852
rect 29596 26012 29652 26068
rect 29932 26236 29988 26292
rect 29260 25004 29316 25060
rect 29372 24780 29428 24836
rect 28588 24668 28644 24724
rect 28364 23938 28420 23940
rect 28364 23886 28366 23938
rect 28366 23886 28418 23938
rect 28418 23886 28420 23938
rect 28364 23884 28420 23886
rect 28252 23772 28308 23828
rect 28140 23660 28196 23716
rect 27692 23212 27748 23268
rect 27692 23042 27748 23044
rect 27692 22990 27694 23042
rect 27694 22990 27746 23042
rect 27746 22990 27748 23042
rect 27692 22988 27748 22990
rect 27244 22876 27300 22932
rect 27468 22146 27524 22148
rect 27468 22094 27470 22146
rect 27470 22094 27522 22146
rect 27522 22094 27524 22146
rect 27468 22092 27524 22094
rect 26572 21644 26628 21700
rect 27580 21698 27636 21700
rect 27580 21646 27582 21698
rect 27582 21646 27634 21698
rect 27634 21646 27636 21698
rect 27580 21644 27636 21646
rect 29596 24780 29652 24836
rect 29484 23548 29540 23604
rect 28700 23042 28756 23044
rect 28700 22990 28702 23042
rect 28702 22990 28754 23042
rect 28754 22990 28756 23042
rect 28700 22988 28756 22990
rect 28588 22594 28644 22596
rect 28588 22542 28590 22594
rect 28590 22542 28642 22594
rect 28642 22542 28644 22594
rect 28588 22540 28644 22542
rect 28476 22428 28532 22484
rect 26908 21586 26964 21588
rect 26908 21534 26910 21586
rect 26910 21534 26962 21586
rect 26962 21534 26964 21586
rect 26908 21532 26964 21534
rect 26684 20972 26740 21028
rect 28476 21644 28532 21700
rect 28364 21586 28420 21588
rect 28364 21534 28366 21586
rect 28366 21534 28418 21586
rect 28418 21534 28420 21586
rect 28364 21532 28420 21534
rect 27692 20802 27748 20804
rect 27692 20750 27694 20802
rect 27694 20750 27746 20802
rect 27746 20750 27748 20802
rect 27692 20748 27748 20750
rect 26572 20076 26628 20132
rect 26684 20018 26740 20020
rect 26684 19966 26686 20018
rect 26686 19966 26738 20018
rect 26738 19966 26740 20018
rect 26684 19964 26740 19966
rect 26460 19628 26516 19684
rect 26572 19740 26628 19796
rect 26236 19122 26292 19124
rect 26236 19070 26238 19122
rect 26238 19070 26290 19122
rect 26290 19070 26292 19122
rect 26236 19068 26292 19070
rect 25788 18396 25844 18452
rect 26348 18284 26404 18340
rect 26348 17836 26404 17892
rect 27244 19852 27300 19908
rect 26796 18396 26852 18452
rect 30380 26178 30436 26180
rect 30380 26126 30382 26178
rect 30382 26126 30434 26178
rect 30434 26126 30436 26178
rect 30380 26124 30436 26126
rect 30716 25564 30772 25620
rect 30828 25506 30884 25508
rect 30828 25454 30830 25506
rect 30830 25454 30882 25506
rect 30882 25454 30884 25506
rect 30828 25452 30884 25454
rect 30268 25394 30324 25396
rect 30268 25342 30270 25394
rect 30270 25342 30322 25394
rect 30322 25342 30324 25394
rect 30268 25340 30324 25342
rect 30492 24834 30548 24836
rect 30492 24782 30494 24834
rect 30494 24782 30546 24834
rect 30546 24782 30548 24834
rect 30492 24780 30548 24782
rect 30380 23938 30436 23940
rect 30380 23886 30382 23938
rect 30382 23886 30434 23938
rect 30434 23886 30436 23938
rect 30380 23884 30436 23886
rect 30492 23826 30548 23828
rect 30492 23774 30494 23826
rect 30494 23774 30546 23826
rect 30546 23774 30548 23826
rect 30492 23772 30548 23774
rect 30268 23660 30324 23716
rect 29708 23324 29764 23380
rect 29036 22876 29092 22932
rect 29484 22594 29540 22596
rect 29484 22542 29486 22594
rect 29486 22542 29538 22594
rect 29538 22542 29540 22594
rect 29484 22540 29540 22542
rect 29932 22988 29988 23044
rect 30156 22482 30212 22484
rect 30156 22430 30158 22482
rect 30158 22430 30210 22482
rect 30210 22430 30212 22482
rect 30156 22428 30212 22430
rect 30044 21756 30100 21812
rect 29260 21698 29316 21700
rect 29260 21646 29262 21698
rect 29262 21646 29314 21698
rect 29314 21646 29316 21698
rect 29260 21644 29316 21646
rect 29708 21586 29764 21588
rect 29708 21534 29710 21586
rect 29710 21534 29762 21586
rect 29762 21534 29764 21586
rect 29708 21532 29764 21534
rect 28924 21196 28980 21252
rect 29260 21026 29316 21028
rect 29260 20974 29262 21026
rect 29262 20974 29314 21026
rect 29314 20974 29316 21026
rect 29260 20972 29316 20974
rect 30156 20748 30212 20804
rect 30604 23548 30660 23604
rect 32060 30882 32116 30884
rect 32060 30830 32062 30882
rect 32062 30830 32114 30882
rect 32114 30830 32116 30882
rect 32060 30828 32116 30830
rect 31948 30716 32004 30772
rect 31276 30210 31332 30212
rect 31276 30158 31278 30210
rect 31278 30158 31330 30210
rect 31330 30158 31332 30210
rect 31276 30156 31332 30158
rect 32396 30994 32452 30996
rect 32396 30942 32398 30994
rect 32398 30942 32450 30994
rect 32450 30942 32452 30994
rect 32396 30940 32452 30942
rect 32284 30380 32340 30436
rect 32396 30156 32452 30212
rect 32060 29650 32116 29652
rect 32060 29598 32062 29650
rect 32062 29598 32114 29650
rect 32114 29598 32116 29650
rect 32060 29596 32116 29598
rect 31388 29538 31444 29540
rect 31388 29486 31390 29538
rect 31390 29486 31442 29538
rect 31442 29486 31444 29538
rect 31388 29484 31444 29486
rect 31724 29260 31780 29316
rect 31500 28754 31556 28756
rect 31500 28702 31502 28754
rect 31502 28702 31554 28754
rect 31554 28702 31556 28754
rect 31500 28700 31556 28702
rect 32172 28588 32228 28644
rect 32508 30044 32564 30100
rect 32732 33516 32788 33572
rect 32732 32732 32788 32788
rect 33180 36652 33236 36708
rect 33404 36482 33460 36484
rect 33404 36430 33406 36482
rect 33406 36430 33458 36482
rect 33458 36430 33460 36482
rect 33404 36428 33460 36430
rect 33292 35420 33348 35476
rect 33740 35698 33796 35700
rect 33740 35646 33742 35698
rect 33742 35646 33794 35698
rect 33794 35646 33796 35698
rect 33740 35644 33796 35646
rect 33628 35532 33684 35588
rect 34076 36876 34132 36932
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35532 36652 35588 36708
rect 36540 36706 36596 36708
rect 36540 36654 36542 36706
rect 36542 36654 36594 36706
rect 36594 36654 36596 36706
rect 36540 36652 36596 36654
rect 34412 36204 34468 36260
rect 35756 36258 35812 36260
rect 35756 36206 35758 36258
rect 35758 36206 35810 36258
rect 35810 36206 35812 36258
rect 35756 36204 35812 36206
rect 33852 35420 33908 35476
rect 34300 35586 34356 35588
rect 34300 35534 34302 35586
rect 34302 35534 34354 35586
rect 34354 35534 34356 35586
rect 34300 35532 34356 35534
rect 33964 34914 34020 34916
rect 33964 34862 33966 34914
rect 33966 34862 34018 34914
rect 34018 34862 34020 34914
rect 33964 34860 34020 34862
rect 34860 35420 34916 35476
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 33628 34130 33684 34132
rect 33628 34078 33630 34130
rect 33630 34078 33682 34130
rect 33682 34078 33684 34130
rect 33628 34076 33684 34078
rect 33068 33516 33124 33572
rect 32956 33292 33012 33348
rect 33740 33628 33796 33684
rect 33628 33458 33684 33460
rect 33628 33406 33630 33458
rect 33630 33406 33682 33458
rect 33682 33406 33684 33458
rect 33628 33404 33684 33406
rect 33628 33180 33684 33236
rect 34188 32732 34244 32788
rect 33404 32620 33460 32676
rect 34076 32674 34132 32676
rect 34076 32622 34078 32674
rect 34078 32622 34130 32674
rect 34130 32622 34132 32674
rect 34076 32620 34132 32622
rect 33180 32508 33236 32564
rect 33628 32562 33684 32564
rect 33628 32510 33630 32562
rect 33630 32510 33682 32562
rect 33682 32510 33684 32562
rect 33628 32508 33684 32510
rect 33180 31948 33236 32004
rect 32508 29484 32564 29540
rect 32508 29036 32564 29092
rect 31724 28476 31780 28532
rect 31164 27804 31220 27860
rect 31500 27746 31556 27748
rect 31500 27694 31502 27746
rect 31502 27694 31554 27746
rect 31554 27694 31556 27746
rect 31500 27692 31556 27694
rect 32508 28530 32564 28532
rect 32508 28478 32510 28530
rect 32510 28478 32562 28530
rect 32562 28478 32564 28530
rect 32508 28476 32564 28478
rect 32396 28028 32452 28084
rect 31948 27858 32004 27860
rect 31948 27806 31950 27858
rect 31950 27806 32002 27858
rect 32002 27806 32004 27858
rect 31948 27804 32004 27806
rect 31948 27132 32004 27188
rect 31164 26290 31220 26292
rect 31164 26238 31166 26290
rect 31166 26238 31218 26290
rect 31218 26238 31220 26290
rect 31164 26236 31220 26238
rect 32172 27692 32228 27748
rect 32284 27580 32340 27636
rect 32844 31164 32900 31220
rect 32620 27804 32676 27860
rect 32732 29148 32788 29204
rect 33068 31500 33124 31556
rect 33292 31106 33348 31108
rect 33292 31054 33294 31106
rect 33294 31054 33346 31106
rect 33346 31054 33348 31106
rect 33292 31052 33348 31054
rect 33068 30828 33124 30884
rect 34188 32562 34244 32564
rect 34188 32510 34190 32562
rect 34190 32510 34242 32562
rect 34242 32510 34244 32562
rect 34188 32508 34244 32510
rect 34076 31554 34132 31556
rect 34076 31502 34078 31554
rect 34078 31502 34130 31554
rect 34130 31502 34132 31554
rect 34076 31500 34132 31502
rect 33404 30268 33460 30324
rect 33516 31388 33572 31444
rect 33180 30156 33236 30212
rect 33740 30994 33796 30996
rect 33740 30942 33742 30994
rect 33742 30942 33794 30994
rect 33794 30942 33796 30994
rect 33740 30940 33796 30942
rect 32956 28924 33012 28980
rect 35084 34076 35140 34132
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35084 33346 35140 33348
rect 35084 33294 35086 33346
rect 35086 33294 35138 33346
rect 35138 33294 35140 33346
rect 35084 33292 35140 33294
rect 34972 33234 35028 33236
rect 34972 33182 34974 33234
rect 34974 33182 35026 33234
rect 35026 33182 35028 33234
rect 34972 33180 35028 33182
rect 34860 30940 34916 30996
rect 34412 29596 34468 29652
rect 34524 30044 34580 30100
rect 33964 29426 34020 29428
rect 33964 29374 33966 29426
rect 33966 29374 34018 29426
rect 34018 29374 34020 29426
rect 33964 29372 34020 29374
rect 33516 29148 33572 29204
rect 33292 28924 33348 28980
rect 33068 28588 33124 28644
rect 33180 28700 33236 28756
rect 32956 28082 33012 28084
rect 32956 28030 32958 28082
rect 32958 28030 33010 28082
rect 33010 28030 33012 28082
rect 32956 28028 33012 28030
rect 33964 28754 34020 28756
rect 33964 28702 33966 28754
rect 33966 28702 34018 28754
rect 34018 28702 34020 28754
rect 33964 28700 34020 28702
rect 33404 28530 33460 28532
rect 33404 28478 33406 28530
rect 33406 28478 33458 28530
rect 33458 28478 33460 28530
rect 33404 28476 33460 28478
rect 32732 27580 32788 27636
rect 33180 27804 33236 27860
rect 31612 26012 31668 26068
rect 31276 25452 31332 25508
rect 31500 25506 31556 25508
rect 31500 25454 31502 25506
rect 31502 25454 31554 25506
rect 31554 25454 31556 25506
rect 31500 25452 31556 25454
rect 31164 25340 31220 25396
rect 31724 24780 31780 24836
rect 31948 26684 32004 26740
rect 32060 25788 32116 25844
rect 31948 25676 32004 25732
rect 31164 23042 31220 23044
rect 31164 22990 31166 23042
rect 31166 22990 31218 23042
rect 31218 22990 31220 23042
rect 31164 22988 31220 22990
rect 31388 22428 31444 22484
rect 31612 22482 31668 22484
rect 31612 22430 31614 22482
rect 31614 22430 31666 22482
rect 31666 22430 31668 22482
rect 31612 22428 31668 22430
rect 30940 21810 30996 21812
rect 30940 21758 30942 21810
rect 30942 21758 30994 21810
rect 30994 21758 30996 21810
rect 30940 21756 30996 21758
rect 30268 21532 30324 21588
rect 28588 20578 28644 20580
rect 28588 20526 28590 20578
rect 28590 20526 28642 20578
rect 28642 20526 28644 20578
rect 28588 20524 28644 20526
rect 29260 20578 29316 20580
rect 29260 20526 29262 20578
rect 29262 20526 29314 20578
rect 29314 20526 29316 20578
rect 29260 20524 29316 20526
rect 30828 21586 30884 21588
rect 30828 21534 30830 21586
rect 30830 21534 30882 21586
rect 30882 21534 30884 21586
rect 30828 21532 30884 21534
rect 30604 20972 30660 21028
rect 29148 20130 29204 20132
rect 29148 20078 29150 20130
rect 29150 20078 29202 20130
rect 29202 20078 29204 20130
rect 29148 20076 29204 20078
rect 29260 19964 29316 20020
rect 30380 20018 30436 20020
rect 30380 19966 30382 20018
rect 30382 19966 30434 20018
rect 30434 19966 30436 20018
rect 30380 19964 30436 19966
rect 25900 17724 25956 17780
rect 25452 17612 25508 17668
rect 25228 17388 25284 17444
rect 25228 17052 25284 17108
rect 26684 17388 26740 17444
rect 26124 16940 26180 16996
rect 25900 16716 25956 16772
rect 24668 15484 24724 15540
rect 23212 14364 23268 14420
rect 22876 12908 22932 12964
rect 22988 12290 23044 12292
rect 22988 12238 22990 12290
rect 22990 12238 23042 12290
rect 23042 12238 23044 12290
rect 22988 12236 23044 12238
rect 22764 12066 22820 12068
rect 22764 12014 22766 12066
rect 22766 12014 22818 12066
rect 22818 12014 22820 12066
rect 22764 12012 22820 12014
rect 22876 11900 22932 11956
rect 22876 10444 22932 10500
rect 22428 9660 22484 9716
rect 23100 11788 23156 11844
rect 23212 9660 23268 9716
rect 22652 7532 22708 7588
rect 22204 6636 22260 6692
rect 22428 6466 22484 6468
rect 22428 6414 22430 6466
rect 22430 6414 22482 6466
rect 22482 6414 22484 6466
rect 22428 6412 22484 6414
rect 21084 3388 21140 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 23100 3554 23156 3556
rect 23100 3502 23102 3554
rect 23102 3502 23154 3554
rect 23154 3502 23156 3554
rect 23100 3500 23156 3502
rect 21756 3442 21812 3444
rect 21756 3390 21758 3442
rect 21758 3390 21810 3442
rect 21810 3390 21812 3442
rect 21756 3388 21812 3390
rect 25788 15538 25844 15540
rect 25788 15486 25790 15538
rect 25790 15486 25842 15538
rect 25842 15486 25844 15538
rect 25788 15484 25844 15486
rect 26012 15932 26068 15988
rect 25340 15260 25396 15316
rect 23996 14364 24052 14420
rect 24108 13970 24164 13972
rect 24108 13918 24110 13970
rect 24110 13918 24162 13970
rect 24162 13918 24164 13970
rect 24108 13916 24164 13918
rect 23772 13804 23828 13860
rect 23772 13132 23828 13188
rect 23884 13634 23940 13636
rect 23884 13582 23886 13634
rect 23886 13582 23938 13634
rect 23938 13582 23940 13634
rect 23884 13580 23940 13582
rect 24332 13580 24388 13636
rect 24220 13468 24276 13524
rect 23660 11900 23716 11956
rect 23772 12236 23828 12292
rect 24780 14476 24836 14532
rect 25228 14140 25284 14196
rect 26572 16940 26628 16996
rect 26796 16940 26852 16996
rect 27356 18338 27412 18340
rect 27356 18286 27358 18338
rect 27358 18286 27410 18338
rect 27410 18286 27412 18338
rect 27356 18284 27412 18286
rect 27580 18284 27636 18340
rect 28476 19234 28532 19236
rect 28476 19182 28478 19234
rect 28478 19182 28530 19234
rect 28530 19182 28532 19234
rect 28476 19180 28532 19182
rect 27020 16716 27076 16772
rect 25676 15148 25732 15204
rect 26684 16044 26740 16100
rect 26348 15820 26404 15876
rect 29932 19794 29988 19796
rect 29932 19742 29934 19794
rect 29934 19742 29986 19794
rect 29986 19742 29988 19794
rect 29932 19740 29988 19742
rect 29708 19628 29764 19684
rect 31052 19628 31108 19684
rect 30156 19180 30212 19236
rect 28028 17388 28084 17444
rect 28476 17276 28532 17332
rect 27804 16940 27860 16996
rect 28476 16940 28532 16996
rect 26908 15874 26964 15876
rect 26908 15822 26910 15874
rect 26910 15822 26962 15874
rect 26962 15822 26964 15874
rect 26908 15820 26964 15822
rect 26908 15260 26964 15316
rect 26124 14812 26180 14868
rect 26236 14588 26292 14644
rect 26124 14530 26180 14532
rect 26124 14478 26126 14530
rect 26126 14478 26178 14530
rect 26178 14478 26180 14530
rect 26124 14476 26180 14478
rect 24780 13020 24836 13076
rect 25452 13634 25508 13636
rect 25452 13582 25454 13634
rect 25454 13582 25506 13634
rect 25506 13582 25508 13634
rect 25452 13580 25508 13582
rect 25228 12796 25284 12852
rect 25340 12908 25396 12964
rect 25228 12178 25284 12180
rect 25228 12126 25230 12178
rect 25230 12126 25282 12178
rect 25282 12126 25284 12178
rect 25228 12124 25284 12126
rect 24556 12012 24612 12068
rect 24444 11282 24500 11284
rect 24444 11230 24446 11282
rect 24446 11230 24498 11282
rect 24498 11230 24500 11282
rect 24444 11228 24500 11230
rect 23772 10668 23828 10724
rect 24332 9826 24388 9828
rect 24332 9774 24334 9826
rect 24334 9774 24386 9826
rect 24386 9774 24388 9826
rect 24332 9772 24388 9774
rect 25452 12796 25508 12852
rect 25452 12124 25508 12180
rect 25004 10332 25060 10388
rect 24780 9884 24836 9940
rect 25228 11228 25284 11284
rect 25340 10722 25396 10724
rect 25340 10670 25342 10722
rect 25342 10670 25394 10722
rect 25394 10670 25396 10722
rect 25340 10668 25396 10670
rect 25116 9996 25172 10052
rect 25452 9772 25508 9828
rect 24780 9266 24836 9268
rect 24780 9214 24782 9266
rect 24782 9214 24834 9266
rect 24834 9214 24836 9266
rect 24780 9212 24836 9214
rect 25228 9602 25284 9604
rect 25228 9550 25230 9602
rect 25230 9550 25282 9602
rect 25282 9550 25284 9602
rect 25228 9548 25284 9550
rect 23436 7586 23492 7588
rect 23436 7534 23438 7586
rect 23438 7534 23490 7586
rect 23490 7534 23492 7586
rect 23436 7532 23492 7534
rect 23772 7586 23828 7588
rect 23772 7534 23774 7586
rect 23774 7534 23826 7586
rect 23826 7534 23828 7586
rect 23772 7532 23828 7534
rect 23772 6690 23828 6692
rect 23772 6638 23774 6690
rect 23774 6638 23826 6690
rect 23826 6638 23828 6690
rect 23772 6636 23828 6638
rect 25116 8034 25172 8036
rect 25116 7982 25118 8034
rect 25118 7982 25170 8034
rect 25170 7982 25172 8034
rect 25116 7980 25172 7982
rect 25340 7532 25396 7588
rect 25676 13020 25732 13076
rect 26012 13186 26068 13188
rect 26012 13134 26014 13186
rect 26014 13134 26066 13186
rect 26066 13134 26068 13186
rect 26012 13132 26068 13134
rect 26236 13132 26292 13188
rect 26348 12908 26404 12964
rect 26012 12684 26068 12740
rect 26572 14364 26628 14420
rect 27244 15986 27300 15988
rect 27244 15934 27246 15986
rect 27246 15934 27298 15986
rect 27298 15934 27300 15986
rect 27244 15932 27300 15934
rect 28140 15820 28196 15876
rect 28700 16882 28756 16884
rect 28700 16830 28702 16882
rect 28702 16830 28754 16882
rect 28754 16830 28756 16882
rect 28700 16828 28756 16830
rect 29148 18338 29204 18340
rect 29148 18286 29150 18338
rect 29150 18286 29202 18338
rect 29202 18286 29204 18338
rect 29148 18284 29204 18286
rect 28588 16098 28644 16100
rect 28588 16046 28590 16098
rect 28590 16046 28642 16098
rect 28642 16046 28644 16098
rect 28588 16044 28644 16046
rect 27132 14700 27188 14756
rect 27244 14588 27300 14644
rect 26796 13916 26852 13972
rect 27020 14476 27076 14532
rect 27580 14700 27636 14756
rect 27916 14754 27972 14756
rect 27916 14702 27918 14754
rect 27918 14702 27970 14754
rect 27970 14702 27972 14754
rect 27916 14700 27972 14702
rect 28028 14588 28084 14644
rect 27020 14306 27076 14308
rect 27020 14254 27022 14306
rect 27022 14254 27074 14306
rect 27074 14254 27076 14306
rect 27020 14252 27076 14254
rect 27916 14252 27972 14308
rect 27356 14140 27412 14196
rect 26684 12684 26740 12740
rect 26684 12012 26740 12068
rect 26460 11900 26516 11956
rect 27020 13580 27076 13636
rect 27020 13356 27076 13412
rect 27244 13356 27300 13412
rect 26908 13186 26964 13188
rect 26908 13134 26910 13186
rect 26910 13134 26962 13186
rect 26962 13134 26964 13186
rect 26908 13132 26964 13134
rect 27132 13074 27188 13076
rect 27132 13022 27134 13074
rect 27134 13022 27186 13074
rect 27186 13022 27188 13074
rect 27132 13020 27188 13022
rect 27132 12684 27188 12740
rect 27020 12066 27076 12068
rect 27020 12014 27022 12066
rect 27022 12014 27074 12066
rect 27074 12014 27076 12066
rect 27020 12012 27076 12014
rect 27244 11900 27300 11956
rect 26908 11452 26964 11508
rect 25900 10332 25956 10388
rect 26460 9884 26516 9940
rect 26572 9826 26628 9828
rect 26572 9774 26574 9826
rect 26574 9774 26626 9826
rect 26626 9774 26628 9826
rect 26572 9772 26628 9774
rect 27468 13020 27524 13076
rect 27580 12850 27636 12852
rect 27580 12798 27582 12850
rect 27582 12798 27634 12850
rect 27634 12798 27636 12850
rect 27580 12796 27636 12798
rect 27804 12962 27860 12964
rect 27804 12910 27806 12962
rect 27806 12910 27858 12962
rect 27858 12910 27860 12962
rect 27804 12908 27860 12910
rect 27692 11506 27748 11508
rect 27692 11454 27694 11506
rect 27694 11454 27746 11506
rect 27746 11454 27748 11506
rect 27692 11452 27748 11454
rect 28252 14418 28308 14420
rect 28252 14366 28254 14418
rect 28254 14366 28306 14418
rect 28306 14366 28308 14418
rect 28252 14364 28308 14366
rect 28364 14306 28420 14308
rect 28364 14254 28366 14306
rect 28366 14254 28418 14306
rect 28418 14254 28420 14306
rect 28364 14252 28420 14254
rect 28140 13858 28196 13860
rect 28140 13806 28142 13858
rect 28142 13806 28194 13858
rect 28194 13806 28196 13858
rect 28140 13804 28196 13806
rect 28028 13580 28084 13636
rect 28140 13356 28196 13412
rect 28028 13132 28084 13188
rect 28140 12738 28196 12740
rect 28140 12686 28142 12738
rect 28142 12686 28194 12738
rect 28194 12686 28196 12738
rect 28140 12684 28196 12686
rect 28028 12572 28084 12628
rect 27132 9996 27188 10052
rect 27020 9772 27076 9828
rect 25900 9324 25956 9380
rect 26796 9548 26852 9604
rect 26012 9212 26068 9268
rect 26460 9154 26516 9156
rect 26460 9102 26462 9154
rect 26462 9102 26514 9154
rect 26514 9102 26516 9154
rect 26460 9100 26516 9102
rect 26908 9100 26964 9156
rect 25900 8034 25956 8036
rect 25900 7982 25902 8034
rect 25902 7982 25954 8034
rect 25954 7982 25956 8034
rect 25900 7980 25956 7982
rect 25788 6636 25844 6692
rect 26012 6412 26068 6468
rect 23548 3554 23604 3556
rect 23548 3502 23550 3554
rect 23550 3502 23602 3554
rect 23602 3502 23604 3554
rect 23548 3500 23604 3502
rect 27132 9436 27188 9492
rect 28364 12962 28420 12964
rect 28364 12910 28366 12962
rect 28366 12910 28418 12962
rect 28418 12910 28420 12962
rect 28364 12908 28420 12910
rect 28252 11676 28308 11732
rect 28252 11116 28308 11172
rect 29372 17778 29428 17780
rect 29372 17726 29374 17778
rect 29374 17726 29426 17778
rect 29426 17726 29428 17778
rect 29372 17724 29428 17726
rect 29260 17612 29316 17668
rect 29708 17666 29764 17668
rect 29708 17614 29710 17666
rect 29710 17614 29762 17666
rect 29762 17614 29764 17666
rect 29708 17612 29764 17614
rect 29260 16044 29316 16100
rect 29260 15874 29316 15876
rect 29260 15822 29262 15874
rect 29262 15822 29314 15874
rect 29314 15822 29316 15874
rect 29260 15820 29316 15822
rect 29820 17276 29876 17332
rect 29820 16940 29876 16996
rect 29596 16098 29652 16100
rect 29596 16046 29598 16098
rect 29598 16046 29650 16098
rect 29650 16046 29652 16098
rect 29596 16044 29652 16046
rect 30044 17724 30100 17780
rect 30716 19234 30772 19236
rect 30716 19182 30718 19234
rect 30718 19182 30770 19234
rect 30770 19182 30772 19234
rect 30716 19180 30772 19182
rect 31500 21756 31556 21812
rect 32508 26460 32564 26516
rect 32844 26124 32900 26180
rect 32060 24444 32116 24500
rect 32508 25282 32564 25284
rect 32508 25230 32510 25282
rect 32510 25230 32562 25282
rect 32562 25230 32564 25282
rect 32508 25228 32564 25230
rect 32396 23884 32452 23940
rect 32172 23324 32228 23380
rect 32284 22258 32340 22260
rect 32284 22206 32286 22258
rect 32286 22206 32338 22258
rect 32338 22206 32340 22258
rect 32284 22204 32340 22206
rect 31836 21362 31892 21364
rect 31836 21310 31838 21362
rect 31838 21310 31890 21362
rect 31890 21310 31892 21362
rect 31836 21308 31892 21310
rect 31724 20860 31780 20916
rect 31276 20524 31332 20580
rect 31500 19964 31556 20020
rect 31276 19794 31332 19796
rect 31276 19742 31278 19794
rect 31278 19742 31330 19794
rect 31330 19742 31332 19794
rect 31276 19740 31332 19742
rect 31052 19122 31108 19124
rect 31052 19070 31054 19122
rect 31054 19070 31106 19122
rect 31106 19070 31108 19122
rect 31052 19068 31108 19070
rect 31164 18844 31220 18900
rect 31500 18844 31556 18900
rect 31724 18338 31780 18340
rect 31724 18286 31726 18338
rect 31726 18286 31778 18338
rect 31778 18286 31780 18338
rect 31724 18284 31780 18286
rect 29932 15932 29988 15988
rect 30268 16044 30324 16100
rect 29820 15596 29876 15652
rect 31388 17612 31444 17668
rect 31388 16828 31444 16884
rect 31052 15986 31108 15988
rect 31052 15934 31054 15986
rect 31054 15934 31106 15986
rect 31106 15934 31108 15986
rect 31052 15932 31108 15934
rect 30604 14812 30660 14868
rect 30716 15820 30772 15876
rect 31164 15372 31220 15428
rect 30828 15202 30884 15204
rect 30828 15150 30830 15202
rect 30830 15150 30882 15202
rect 30882 15150 30884 15202
rect 30828 15148 30884 15150
rect 31052 15314 31108 15316
rect 31052 15262 31054 15314
rect 31054 15262 31106 15314
rect 31106 15262 31108 15314
rect 31052 15260 31108 15262
rect 29708 14530 29764 14532
rect 29708 14478 29710 14530
rect 29710 14478 29762 14530
rect 29762 14478 29764 14530
rect 29708 14476 29764 14478
rect 30716 14588 30772 14644
rect 31052 15036 31108 15092
rect 28924 14364 28980 14420
rect 29148 13804 29204 13860
rect 29596 13356 29652 13412
rect 30604 13804 30660 13860
rect 30380 13468 30436 13524
rect 28812 12572 28868 12628
rect 29372 12572 29428 12628
rect 28924 12290 28980 12292
rect 28924 12238 28926 12290
rect 28926 12238 28978 12290
rect 28978 12238 28980 12290
rect 28924 12236 28980 12238
rect 29708 13132 29764 13188
rect 28476 12178 28532 12180
rect 28476 12126 28478 12178
rect 28478 12126 28530 12178
rect 28530 12126 28532 12178
rect 28476 12124 28532 12126
rect 28476 11394 28532 11396
rect 28476 11342 28478 11394
rect 28478 11342 28530 11394
rect 28530 11342 28532 11394
rect 28476 11340 28532 11342
rect 28364 10668 28420 10724
rect 27580 9996 27636 10052
rect 28476 9100 28532 9156
rect 28924 9212 28980 9268
rect 29596 12124 29652 12180
rect 29484 11676 29540 11732
rect 29260 11170 29316 11172
rect 29260 11118 29262 11170
rect 29262 11118 29314 11170
rect 29314 11118 29316 11170
rect 29260 11116 29316 11118
rect 30492 13132 30548 13188
rect 29932 12236 29988 12292
rect 29820 11340 29876 11396
rect 30044 12178 30100 12180
rect 30044 12126 30046 12178
rect 30046 12126 30098 12178
rect 30098 12126 30100 12178
rect 30044 12124 30100 12126
rect 30940 14252 30996 14308
rect 30940 13692 30996 13748
rect 31052 14476 31108 14532
rect 31164 13468 31220 13524
rect 30828 13132 30884 13188
rect 30716 13020 30772 13076
rect 30604 12572 30660 12628
rect 30604 12290 30660 12292
rect 30604 12238 30606 12290
rect 30606 12238 30658 12290
rect 30658 12238 30660 12290
rect 30604 12236 30660 12238
rect 30716 12124 30772 12180
rect 30828 12012 30884 12068
rect 30380 11340 30436 11396
rect 30044 9996 30100 10052
rect 30940 11452 30996 11508
rect 30604 11228 30660 11284
rect 30604 10332 30660 10388
rect 29260 9772 29316 9828
rect 30156 9772 30212 9828
rect 29260 9324 29316 9380
rect 30044 9602 30100 9604
rect 30044 9550 30046 9602
rect 30046 9550 30098 9602
rect 30098 9550 30100 9602
rect 30044 9548 30100 9550
rect 29372 9436 29428 9492
rect 29596 9324 29652 9380
rect 28140 8204 28196 8260
rect 27468 8146 27524 8148
rect 27468 8094 27470 8146
rect 27470 8094 27522 8146
rect 27522 8094 27524 8146
rect 27468 8092 27524 8094
rect 28028 8146 28084 8148
rect 28028 8094 28030 8146
rect 28030 8094 28082 8146
rect 28082 8094 28084 8146
rect 28028 8092 28084 8094
rect 26796 6524 26852 6580
rect 29148 8258 29204 8260
rect 29148 8206 29150 8258
rect 29150 8206 29202 8258
rect 29202 8206 29204 8258
rect 29148 8204 29204 8206
rect 29372 9100 29428 9156
rect 29372 8316 29428 8372
rect 29708 8764 29764 8820
rect 31724 16604 31780 16660
rect 31612 16044 31668 16100
rect 31500 15202 31556 15204
rect 31500 15150 31502 15202
rect 31502 15150 31554 15202
rect 31554 15150 31556 15202
rect 31500 15148 31556 15150
rect 32060 20524 32116 20580
rect 31948 20018 32004 20020
rect 31948 19966 31950 20018
rect 31950 19966 32002 20018
rect 32002 19966 32004 20018
rect 31948 19964 32004 19966
rect 34300 28642 34356 28644
rect 34300 28590 34302 28642
rect 34302 28590 34354 28642
rect 34354 28590 34356 28642
rect 34300 28588 34356 28590
rect 34748 29036 34804 29092
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 39564 31666 39620 31668
rect 39564 31614 39566 31666
rect 39566 31614 39618 31666
rect 39618 31614 39620 31666
rect 39564 31612 39620 31614
rect 40012 31612 40068 31668
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35420 30380 35476 30436
rect 35196 29426 35252 29428
rect 35196 29374 35198 29426
rect 35198 29374 35250 29426
rect 35250 29374 35252 29426
rect 35196 29372 35252 29374
rect 35644 30268 35700 30324
rect 39900 31388 39956 31444
rect 40236 30994 40292 30996
rect 40236 30942 40238 30994
rect 40238 30942 40290 30994
rect 40290 30942 40292 30994
rect 40236 30940 40292 30942
rect 39228 30268 39284 30324
rect 37100 29596 37156 29652
rect 34972 29314 35028 29316
rect 34972 29262 34974 29314
rect 34974 29262 35026 29314
rect 35026 29262 35028 29314
rect 34972 29260 35028 29262
rect 35868 29314 35924 29316
rect 35868 29262 35870 29314
rect 35870 29262 35922 29314
rect 35922 29262 35924 29314
rect 35868 29260 35924 29262
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35532 28812 35588 28868
rect 35420 28700 35476 28756
rect 36316 28642 36372 28644
rect 36316 28590 36318 28642
rect 36318 28590 36370 28642
rect 36370 28590 36372 28642
rect 36316 28588 36372 28590
rect 37100 28642 37156 28644
rect 37100 28590 37102 28642
rect 37102 28590 37154 28642
rect 37154 28590 37156 28642
rect 37100 28588 37156 28590
rect 37436 29372 37492 29428
rect 39004 29426 39060 29428
rect 39004 29374 39006 29426
rect 39006 29374 39058 29426
rect 39058 29374 39060 29426
rect 39004 29372 39060 29374
rect 37436 28700 37492 28756
rect 34636 28476 34692 28532
rect 34412 28364 34468 28420
rect 33740 27858 33796 27860
rect 33740 27806 33742 27858
rect 33742 27806 33794 27858
rect 33794 27806 33796 27858
rect 33740 27804 33796 27806
rect 33516 27244 33572 27300
rect 36092 28418 36148 28420
rect 36092 28366 36094 28418
rect 36094 28366 36146 28418
rect 36146 28366 36148 28418
rect 36092 28364 36148 28366
rect 39900 29148 39956 29204
rect 37548 28642 37604 28644
rect 37548 28590 37550 28642
rect 37550 28590 37602 28642
rect 37602 28590 37604 28642
rect 37548 28588 37604 28590
rect 40124 28924 40180 28980
rect 39676 28252 39732 28308
rect 40236 28252 40292 28308
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 33404 27186 33460 27188
rect 33404 27134 33406 27186
rect 33406 27134 33458 27186
rect 33458 27134 33460 27186
rect 33404 27132 33460 27134
rect 34748 27244 34804 27300
rect 33404 26514 33460 26516
rect 33404 26462 33406 26514
rect 33406 26462 33458 26514
rect 33458 26462 33460 26514
rect 33404 26460 33460 26462
rect 32956 25676 33012 25732
rect 34412 26684 34468 26740
rect 33964 26290 34020 26292
rect 33964 26238 33966 26290
rect 33966 26238 34018 26290
rect 34018 26238 34020 26290
rect 33964 26236 34020 26238
rect 36540 26236 36596 26292
rect 33292 26124 33348 26180
rect 33516 26066 33572 26068
rect 33516 26014 33518 26066
rect 33518 26014 33570 26066
rect 33570 26014 33572 26066
rect 33516 26012 33572 26014
rect 33292 25788 33348 25844
rect 33068 24834 33124 24836
rect 33068 24782 33070 24834
rect 33070 24782 33122 24834
rect 33122 24782 33124 24834
rect 33068 24780 33124 24782
rect 33180 24668 33236 24724
rect 33068 23938 33124 23940
rect 33068 23886 33070 23938
rect 33070 23886 33122 23938
rect 33122 23886 33124 23938
rect 33068 23884 33124 23886
rect 33516 24444 33572 24500
rect 33292 23378 33348 23380
rect 33292 23326 33294 23378
rect 33294 23326 33346 23378
rect 33346 23326 33348 23378
rect 33292 23324 33348 23326
rect 32844 22428 32900 22484
rect 32956 22370 33012 22372
rect 32956 22318 32958 22370
rect 32958 22318 33010 22370
rect 33010 22318 33012 22370
rect 32956 22316 33012 22318
rect 35308 26012 35364 26068
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34860 25676 34916 25732
rect 35756 25676 35812 25732
rect 34636 24780 34692 24836
rect 34188 24668 34244 24724
rect 34412 24610 34468 24612
rect 34412 24558 34414 24610
rect 34414 24558 34466 24610
rect 34466 24558 34468 24610
rect 34412 24556 34468 24558
rect 34300 23884 34356 23940
rect 39004 26290 39060 26292
rect 39004 26238 39006 26290
rect 39006 26238 39058 26290
rect 39058 26238 39060 26290
rect 39004 26236 39060 26238
rect 36540 25730 36596 25732
rect 36540 25678 36542 25730
rect 36542 25678 36594 25730
rect 36594 25678 36596 25730
rect 36540 25676 36596 25678
rect 40124 25564 40180 25620
rect 39004 25506 39060 25508
rect 39004 25454 39006 25506
rect 39006 25454 39058 25506
rect 39058 25454 39060 25506
rect 39004 25452 39060 25454
rect 35756 25228 35812 25284
rect 39788 24892 39844 24948
rect 36204 24834 36260 24836
rect 36204 24782 36206 24834
rect 36206 24782 36258 24834
rect 36258 24782 36260 24834
rect 36204 24780 36260 24782
rect 36316 24722 36372 24724
rect 36316 24670 36318 24722
rect 36318 24670 36370 24722
rect 36370 24670 36372 24722
rect 36316 24668 36372 24670
rect 35644 24556 35700 24612
rect 35420 24444 35476 24500
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 33516 22316 33572 22372
rect 33404 22258 33460 22260
rect 33404 22206 33406 22258
rect 33406 22206 33458 22258
rect 33458 22206 33460 22258
rect 33404 22204 33460 22206
rect 35420 23938 35476 23940
rect 35420 23886 35422 23938
rect 35422 23886 35474 23938
rect 35474 23886 35476 23938
rect 35420 23884 35476 23886
rect 35868 23938 35924 23940
rect 35868 23886 35870 23938
rect 35870 23886 35922 23938
rect 35922 23886 35924 23938
rect 35868 23884 35924 23886
rect 39004 23938 39060 23940
rect 39004 23886 39006 23938
rect 39006 23886 39058 23938
rect 39058 23886 39060 23938
rect 39004 23884 39060 23886
rect 36764 23548 36820 23604
rect 38332 23548 38388 23604
rect 34076 23266 34132 23268
rect 34076 23214 34078 23266
rect 34078 23214 34130 23266
rect 34130 23214 34132 23266
rect 34076 23212 34132 23214
rect 34636 23266 34692 23268
rect 34636 23214 34638 23266
rect 34638 23214 34690 23266
rect 34690 23214 34692 23266
rect 34636 23212 34692 23214
rect 33852 22258 33908 22260
rect 33852 22206 33854 22258
rect 33854 22206 33906 22258
rect 33906 22206 33908 22258
rect 33852 22204 33908 22206
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35084 22428 35140 22484
rect 34972 22370 35028 22372
rect 34972 22318 34974 22370
rect 34974 22318 35026 22370
rect 35026 22318 35028 22370
rect 34972 22316 35028 22318
rect 33180 21980 33236 22036
rect 33292 21868 33348 21924
rect 32732 21756 32788 21812
rect 32508 21586 32564 21588
rect 32508 21534 32510 21586
rect 32510 21534 32562 21586
rect 32562 21534 32564 21586
rect 32508 21532 32564 21534
rect 33292 21362 33348 21364
rect 33292 21310 33294 21362
rect 33294 21310 33346 21362
rect 33346 21310 33348 21362
rect 33292 21308 33348 21310
rect 33740 21810 33796 21812
rect 33740 21758 33742 21810
rect 33742 21758 33794 21810
rect 33794 21758 33796 21810
rect 33740 21756 33796 21758
rect 33628 21644 33684 21700
rect 33852 21698 33908 21700
rect 33852 21646 33854 21698
rect 33854 21646 33906 21698
rect 33906 21646 33908 21698
rect 33852 21644 33908 21646
rect 33628 20914 33684 20916
rect 33628 20862 33630 20914
rect 33630 20862 33682 20914
rect 33682 20862 33684 20914
rect 33628 20860 33684 20862
rect 32844 20802 32900 20804
rect 32844 20750 32846 20802
rect 32846 20750 32898 20802
rect 32898 20750 32900 20802
rect 32844 20748 32900 20750
rect 33964 21586 34020 21588
rect 33964 21534 33966 21586
rect 33966 21534 34018 21586
rect 34018 21534 34020 21586
rect 33964 21532 34020 21534
rect 33740 20636 33796 20692
rect 32284 19964 32340 20020
rect 32620 20578 32676 20580
rect 32620 20526 32622 20578
rect 32622 20526 32674 20578
rect 32674 20526 32676 20578
rect 32620 20524 32676 20526
rect 34636 21644 34692 21700
rect 34412 20860 34468 20916
rect 32508 19740 32564 19796
rect 32620 19122 32676 19124
rect 32620 19070 32622 19122
rect 32622 19070 32674 19122
rect 32674 19070 32676 19122
rect 32620 19068 32676 19070
rect 32732 18844 32788 18900
rect 32172 18338 32228 18340
rect 32172 18286 32174 18338
rect 32174 18286 32226 18338
rect 32226 18286 32228 18338
rect 32172 18284 32228 18286
rect 33628 19516 33684 19572
rect 33516 18844 33572 18900
rect 33740 18284 33796 18340
rect 35868 22482 35924 22484
rect 35868 22430 35870 22482
rect 35870 22430 35922 22482
rect 35922 22430 35924 22482
rect 35868 22428 35924 22430
rect 35420 22258 35476 22260
rect 35420 22206 35422 22258
rect 35422 22206 35474 22258
rect 35474 22206 35476 22258
rect 35420 22204 35476 22206
rect 40012 23548 40068 23604
rect 38556 23042 38612 23044
rect 38556 22990 38558 23042
rect 38558 22990 38610 23042
rect 38610 22990 38612 23042
rect 38556 22988 38612 22990
rect 35084 21308 35140 21364
rect 37996 21532 38052 21588
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35420 21026 35476 21028
rect 35420 20974 35422 21026
rect 35422 20974 35474 21026
rect 35474 20974 35476 21026
rect 35420 20972 35476 20974
rect 37996 20972 38052 21028
rect 35532 20914 35588 20916
rect 35532 20862 35534 20914
rect 35534 20862 35586 20914
rect 35586 20862 35588 20914
rect 35532 20860 35588 20862
rect 35084 20802 35140 20804
rect 35084 20750 35086 20802
rect 35086 20750 35138 20802
rect 35138 20750 35140 20802
rect 35084 20748 35140 20750
rect 35196 20636 35252 20692
rect 34524 20524 34580 20580
rect 34972 20524 35028 20580
rect 34188 20076 34244 20132
rect 36092 20578 36148 20580
rect 36092 20526 36094 20578
rect 36094 20526 36146 20578
rect 36146 20526 36148 20578
rect 36092 20524 36148 20526
rect 33852 18172 33908 18228
rect 34076 19068 34132 19124
rect 34748 18284 34804 18340
rect 34524 18226 34580 18228
rect 34524 18174 34526 18226
rect 34526 18174 34578 18226
rect 34578 18174 34580 18226
rect 34524 18172 34580 18174
rect 32844 17442 32900 17444
rect 32844 17390 32846 17442
rect 32846 17390 32898 17442
rect 32898 17390 32900 17442
rect 32844 17388 32900 17390
rect 32060 17052 32116 17108
rect 32396 15874 32452 15876
rect 32396 15822 32398 15874
rect 32398 15822 32450 15874
rect 32450 15822 32452 15874
rect 32396 15820 32452 15822
rect 32060 15708 32116 15764
rect 33292 16994 33348 16996
rect 33292 16942 33294 16994
rect 33294 16942 33346 16994
rect 33346 16942 33348 16994
rect 33292 16940 33348 16942
rect 33180 16658 33236 16660
rect 33180 16606 33182 16658
rect 33182 16606 33234 16658
rect 33234 16606 33236 16658
rect 33180 16604 33236 16606
rect 33292 16156 33348 16212
rect 33292 15986 33348 15988
rect 33292 15934 33294 15986
rect 33294 15934 33346 15986
rect 33346 15934 33348 15986
rect 33292 15932 33348 15934
rect 32284 15596 32340 15652
rect 32060 15260 32116 15316
rect 32172 15484 32228 15540
rect 31500 14812 31556 14868
rect 32620 15260 32676 15316
rect 32956 15708 33012 15764
rect 33404 15874 33460 15876
rect 33404 15822 33406 15874
rect 33406 15822 33458 15874
rect 33458 15822 33460 15874
rect 33404 15820 33460 15822
rect 33628 16882 33684 16884
rect 33628 16830 33630 16882
rect 33630 16830 33682 16882
rect 33682 16830 33684 16882
rect 33628 16828 33684 16830
rect 34188 16940 34244 16996
rect 32620 14924 32676 14980
rect 32508 13858 32564 13860
rect 32508 13806 32510 13858
rect 32510 13806 32562 13858
rect 32562 13806 32564 13858
rect 32508 13804 32564 13806
rect 31612 13746 31668 13748
rect 31612 13694 31614 13746
rect 31614 13694 31666 13746
rect 31666 13694 31668 13746
rect 31612 13692 31668 13694
rect 32060 13580 32116 13636
rect 32284 13746 32340 13748
rect 32284 13694 32286 13746
rect 32286 13694 32338 13746
rect 32338 13694 32340 13746
rect 32284 13692 32340 13694
rect 31164 11394 31220 11396
rect 31164 11342 31166 11394
rect 31166 11342 31218 11394
rect 31218 11342 31220 11394
rect 31164 11340 31220 11342
rect 31052 11282 31108 11284
rect 31052 11230 31054 11282
rect 31054 11230 31106 11282
rect 31106 11230 31108 11282
rect 31052 11228 31108 11230
rect 31276 11282 31332 11284
rect 31276 11230 31278 11282
rect 31278 11230 31330 11282
rect 31330 11230 31332 11282
rect 31276 11228 31332 11230
rect 30940 10780 30996 10836
rect 31276 10834 31332 10836
rect 31276 10782 31278 10834
rect 31278 10782 31330 10834
rect 31330 10782 31332 10834
rect 31276 10780 31332 10782
rect 30716 9660 30772 9716
rect 30380 9266 30436 9268
rect 30380 9214 30382 9266
rect 30382 9214 30434 9266
rect 30434 9214 30436 9266
rect 30380 9212 30436 9214
rect 30828 9602 30884 9604
rect 30828 9550 30830 9602
rect 30830 9550 30882 9602
rect 30882 9550 30884 9602
rect 30828 9548 30884 9550
rect 32732 13692 32788 13748
rect 33964 15820 34020 15876
rect 34636 17778 34692 17780
rect 34636 17726 34638 17778
rect 34638 17726 34690 17778
rect 34690 17726 34692 17778
rect 34636 17724 34692 17726
rect 34524 17442 34580 17444
rect 34524 17390 34526 17442
rect 34526 17390 34578 17442
rect 34578 17390 34580 17442
rect 34524 17388 34580 17390
rect 34636 16322 34692 16324
rect 34636 16270 34638 16322
rect 34638 16270 34690 16322
rect 34690 16270 34692 16322
rect 34636 16268 34692 16270
rect 34524 15986 34580 15988
rect 34524 15934 34526 15986
rect 34526 15934 34578 15986
rect 34578 15934 34580 15986
rect 34524 15932 34580 15934
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35532 19404 35588 19460
rect 39116 21532 39172 21588
rect 39004 20412 39060 20468
rect 38444 20130 38500 20132
rect 38444 20078 38446 20130
rect 38446 20078 38498 20130
rect 38498 20078 38500 20130
rect 38444 20076 38500 20078
rect 40236 22876 40292 22932
rect 40012 22204 40068 22260
rect 39900 22092 39956 22148
rect 39564 21532 39620 21588
rect 40124 20860 40180 20916
rect 39676 20188 39732 20244
rect 39228 20076 39284 20132
rect 35532 18338 35588 18340
rect 35532 18286 35534 18338
rect 35534 18286 35586 18338
rect 35586 18286 35588 18338
rect 35532 18284 35588 18286
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35980 17778 36036 17780
rect 35980 17726 35982 17778
rect 35982 17726 36034 17778
rect 36034 17726 36036 17778
rect 35980 17724 36036 17726
rect 34972 17500 35028 17556
rect 35532 17554 35588 17556
rect 35532 17502 35534 17554
rect 35534 17502 35586 17554
rect 35586 17502 35588 17554
rect 35532 17500 35588 17502
rect 34860 16828 34916 16884
rect 34412 15708 34468 15764
rect 34860 15708 34916 15764
rect 33740 15372 33796 15428
rect 33180 15036 33236 15092
rect 32956 14418 33012 14420
rect 32956 14366 32958 14418
rect 32958 14366 33010 14418
rect 33010 14366 33012 14418
rect 32956 14364 33012 14366
rect 33068 13916 33124 13972
rect 33628 15314 33684 15316
rect 33628 15262 33630 15314
rect 33630 15262 33682 15314
rect 33682 15262 33684 15314
rect 33628 15260 33684 15262
rect 33292 14924 33348 14980
rect 32844 13580 32900 13636
rect 32732 13186 32788 13188
rect 32732 13134 32734 13186
rect 32734 13134 32786 13186
rect 32786 13134 32788 13186
rect 32732 13132 32788 13134
rect 34188 14364 34244 14420
rect 34188 13916 34244 13972
rect 34636 15260 34692 15316
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35532 16210 35588 16212
rect 35532 16158 35534 16210
rect 35534 16158 35586 16210
rect 35586 16158 35588 16210
rect 35532 16156 35588 16158
rect 37212 16994 37268 16996
rect 37212 16942 37214 16994
rect 37214 16942 37266 16994
rect 37266 16942 37268 16994
rect 37212 16940 37268 16942
rect 35084 15874 35140 15876
rect 35084 15822 35086 15874
rect 35086 15822 35138 15874
rect 35138 15822 35140 15874
rect 35084 15820 35140 15822
rect 35532 15820 35588 15876
rect 34748 15090 34804 15092
rect 34748 15038 34750 15090
rect 34750 15038 34802 15090
rect 34802 15038 34804 15090
rect 34748 15036 34804 15038
rect 34636 14924 34692 14980
rect 33516 13132 33572 13188
rect 33068 12796 33124 12852
rect 30940 9436 30996 9492
rect 30268 8764 30324 8820
rect 30604 8370 30660 8372
rect 30604 8318 30606 8370
rect 30606 8318 30658 8370
rect 30658 8318 30660 8370
rect 30604 8316 30660 8318
rect 28700 7586 28756 7588
rect 28700 7534 28702 7586
rect 28702 7534 28754 7586
rect 28754 7534 28756 7586
rect 28700 7532 28756 7534
rect 33628 12348 33684 12404
rect 33740 12290 33796 12292
rect 33740 12238 33742 12290
rect 33742 12238 33794 12290
rect 33794 12238 33796 12290
rect 33740 12236 33796 12238
rect 32060 11900 32116 11956
rect 31836 11340 31892 11396
rect 30940 8316 30996 8372
rect 31164 8370 31220 8372
rect 31164 8318 31166 8370
rect 31166 8318 31218 8370
rect 31218 8318 31220 8370
rect 31164 8316 31220 8318
rect 31612 10722 31668 10724
rect 31612 10670 31614 10722
rect 31614 10670 31666 10722
rect 31666 10670 31668 10722
rect 31612 10668 31668 10670
rect 31500 9660 31556 9716
rect 31388 9436 31444 9492
rect 31500 9154 31556 9156
rect 31500 9102 31502 9154
rect 31502 9102 31554 9154
rect 31554 9102 31556 9154
rect 31500 9100 31556 9102
rect 31612 9042 31668 9044
rect 31612 8990 31614 9042
rect 31614 8990 31666 9042
rect 31666 8990 31668 9042
rect 31612 8988 31668 8990
rect 34524 13634 34580 13636
rect 34524 13582 34526 13634
rect 34526 13582 34578 13634
rect 34578 13582 34580 13634
rect 34524 13580 34580 13582
rect 34076 13468 34132 13524
rect 34188 13132 34244 13188
rect 34524 12796 34580 12852
rect 34188 12684 34244 12740
rect 33964 11900 34020 11956
rect 34076 12236 34132 12292
rect 34076 11788 34132 11844
rect 33404 11452 33460 11508
rect 35756 15036 35812 15092
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34860 14252 34916 14308
rect 34748 12962 34804 12964
rect 34748 12910 34750 12962
rect 34750 12910 34802 12962
rect 34802 12910 34804 12962
rect 34748 12908 34804 12910
rect 33740 11340 33796 11396
rect 32284 10332 32340 10388
rect 32060 9996 32116 10052
rect 32284 9714 32340 9716
rect 32284 9662 32286 9714
rect 32286 9662 32338 9714
rect 32338 9662 32340 9714
rect 32284 9660 32340 9662
rect 31948 9548 32004 9604
rect 32844 9660 32900 9716
rect 33964 11228 34020 11284
rect 34300 11170 34356 11172
rect 34300 11118 34302 11170
rect 34302 11118 34354 11170
rect 34354 11118 34356 11170
rect 34300 11116 34356 11118
rect 34636 12684 34692 12740
rect 34524 12402 34580 12404
rect 34524 12350 34526 12402
rect 34526 12350 34578 12402
rect 34578 12350 34580 12402
rect 34524 12348 34580 12350
rect 34748 12178 34804 12180
rect 34748 12126 34750 12178
rect 34750 12126 34802 12178
rect 34802 12126 34804 12178
rect 34748 12124 34804 12126
rect 34636 12066 34692 12068
rect 34636 12014 34638 12066
rect 34638 12014 34690 12066
rect 34690 12014 34692 12066
rect 34636 12012 34692 12014
rect 34524 11394 34580 11396
rect 34524 11342 34526 11394
rect 34526 11342 34578 11394
rect 34578 11342 34580 11394
rect 34524 11340 34580 11342
rect 34300 10332 34356 10388
rect 34636 10050 34692 10052
rect 34636 9998 34638 10050
rect 34638 9998 34690 10050
rect 34690 9998 34692 10050
rect 34636 9996 34692 9998
rect 33516 9884 33572 9940
rect 32284 9212 32340 9268
rect 32060 9042 32116 9044
rect 32060 8990 32062 9042
rect 32062 8990 32114 9042
rect 32114 8990 32116 9042
rect 32060 8988 32116 8990
rect 31836 8876 31892 8932
rect 31500 8818 31556 8820
rect 31500 8766 31502 8818
rect 31502 8766 31554 8818
rect 31554 8766 31556 8818
rect 31500 8764 31556 8766
rect 32620 9042 32676 9044
rect 32620 8990 32622 9042
rect 32622 8990 32674 9042
rect 32674 8990 32676 9042
rect 32620 8988 32676 8990
rect 33068 8876 33124 8932
rect 31724 8370 31780 8372
rect 31724 8318 31726 8370
rect 31726 8318 31778 8370
rect 31778 8318 31780 8370
rect 31724 8316 31780 8318
rect 31276 8204 31332 8260
rect 32620 8258 32676 8260
rect 32620 8206 32622 8258
rect 32622 8206 32674 8258
rect 32674 8206 32676 8258
rect 32620 8204 32676 8206
rect 33068 8204 33124 8260
rect 31948 8092 32004 8148
rect 31836 7586 31892 7588
rect 31836 7534 31838 7586
rect 31838 7534 31890 7586
rect 31890 7534 31892 7586
rect 31836 7532 31892 7534
rect 33964 9772 34020 9828
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35644 13692 35700 13748
rect 35532 13132 35588 13188
rect 34972 12850 35028 12852
rect 34972 12798 34974 12850
rect 34974 12798 35026 12850
rect 35026 12798 35028 12850
rect 34972 12796 35028 12798
rect 36092 14306 36148 14308
rect 36092 14254 36094 14306
rect 36094 14254 36146 14306
rect 36146 14254 36148 14306
rect 36092 14252 36148 14254
rect 40236 20188 40292 20244
rect 40012 19516 40068 19572
rect 39900 19292 39956 19348
rect 39900 19010 39956 19012
rect 39900 18958 39902 19010
rect 39902 18958 39954 19010
rect 39954 18958 39956 19010
rect 39900 18956 39956 18958
rect 39676 18844 39732 18900
rect 40236 18844 40292 18900
rect 39004 16268 39060 16324
rect 39004 16098 39060 16100
rect 39004 16046 39006 16098
rect 39006 16046 39058 16098
rect 39058 16046 39060 16098
rect 39004 16044 39060 16046
rect 40012 16828 40068 16884
rect 39788 16156 39844 16212
rect 39116 15484 39172 15540
rect 39228 15708 39284 15764
rect 39004 14700 39060 14756
rect 40124 15484 40180 15540
rect 39788 14812 39844 14868
rect 40236 14140 40292 14196
rect 38556 13970 38612 13972
rect 38556 13918 38558 13970
rect 38558 13918 38610 13970
rect 38610 13918 38612 13970
rect 38556 13916 38612 13918
rect 38668 13692 38724 13748
rect 35980 12962 36036 12964
rect 35980 12910 35982 12962
rect 35982 12910 36034 12962
rect 36034 12910 36036 12962
rect 35980 12908 36036 12910
rect 34972 12290 35028 12292
rect 34972 12238 34974 12290
rect 34974 12238 35026 12290
rect 35026 12238 35028 12290
rect 34972 12236 35028 12238
rect 36204 12738 36260 12740
rect 36204 12686 36206 12738
rect 36206 12686 36258 12738
rect 36258 12686 36260 12738
rect 36204 12684 36260 12686
rect 35980 12348 36036 12404
rect 35196 11900 35252 11956
rect 35532 11900 35588 11956
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34972 11340 35028 11396
rect 35980 11900 36036 11956
rect 35084 11282 35140 11284
rect 35084 11230 35086 11282
rect 35086 11230 35138 11282
rect 35138 11230 35140 11282
rect 35084 11228 35140 11230
rect 33852 9154 33908 9156
rect 33852 9102 33854 9154
rect 33854 9102 33906 9154
rect 33906 9102 33908 9154
rect 33852 9100 33908 9102
rect 34188 9660 34244 9716
rect 34076 9266 34132 9268
rect 34076 9214 34078 9266
rect 34078 9214 34130 9266
rect 34130 9214 34132 9266
rect 34076 9212 34132 9214
rect 34636 9714 34692 9716
rect 34636 9662 34638 9714
rect 34638 9662 34690 9714
rect 34690 9662 34692 9714
rect 34636 9660 34692 9662
rect 34748 9548 34804 9604
rect 35308 10332 35364 10388
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35532 9772 35588 9828
rect 36092 11282 36148 11284
rect 36092 11230 36094 11282
rect 36094 11230 36146 11282
rect 36146 11230 36148 11282
rect 36092 11228 36148 11230
rect 37212 11282 37268 11284
rect 37212 11230 37214 11282
rect 37214 11230 37266 11282
rect 37266 11230 37268 11282
rect 37212 11228 37268 11230
rect 40012 13468 40068 13524
rect 39452 12850 39508 12852
rect 39452 12798 39454 12850
rect 39454 12798 39506 12850
rect 39506 12798 39508 12850
rect 39452 12796 39508 12798
rect 40236 12850 40292 12852
rect 40236 12798 40238 12850
rect 40238 12798 40290 12850
rect 40290 12798 40292 12850
rect 40236 12796 40292 12798
rect 39676 12348 39732 12404
rect 37660 10668 37716 10724
rect 36204 9548 36260 9604
rect 36316 9660 36372 9716
rect 35084 9266 35140 9268
rect 35084 9214 35086 9266
rect 35086 9214 35138 9266
rect 35138 9214 35140 9266
rect 35084 9212 35140 9214
rect 33964 8988 34020 9044
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 32396 7586 32452 7588
rect 32396 7534 32398 7586
rect 32398 7534 32450 7586
rect 32450 7534 32452 7586
rect 32396 7532 32452 7534
rect 35420 7586 35476 7588
rect 35420 7534 35422 7586
rect 35422 7534 35474 7586
rect 35474 7534 35476 7586
rect 35420 7532 35476 7534
rect 35868 7586 35924 7588
rect 35868 7534 35870 7586
rect 35870 7534 35922 7586
rect 35922 7534 35924 7586
rect 35868 7532 35924 7534
rect 38668 10722 38724 10724
rect 38668 10670 38670 10722
rect 38670 10670 38722 10722
rect 38722 10670 38724 10722
rect 38668 10668 38724 10670
rect 39116 10722 39172 10724
rect 39116 10670 39118 10722
rect 39118 10670 39170 10722
rect 39170 10670 39172 10722
rect 39116 10668 39172 10670
rect 37660 7532 37716 7588
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 28364 6690 28420 6692
rect 28364 6638 28366 6690
rect 28366 6638 28418 6690
rect 28418 6638 28420 6690
rect 28364 6636 28420 6638
rect 31724 6636 31780 6692
rect 27804 6524 27860 6580
rect 27916 6466 27972 6468
rect 27916 6414 27918 6466
rect 27918 6414 27970 6466
rect 27970 6414 27972 6466
rect 27916 6412 27972 6414
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
<< metal3 >>
rect 26226 38556 26236 38612
rect 26292 38556 28812 38612
rect 28868 38556 28878 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 12674 38332 12684 38388
rect 12740 38332 16716 38388
rect 16772 38332 17500 38388
rect 17556 38332 17566 38388
rect 14802 38220 14812 38276
rect 14868 38220 15484 38276
rect 15540 38220 15550 38276
rect 18162 38220 18172 38276
rect 18228 38220 19516 38276
rect 19572 38220 19582 38276
rect 28914 38220 28924 38276
rect 28980 38220 30380 38276
rect 30436 38220 30446 38276
rect 10994 37996 11004 38052
rect 11060 37996 11676 38052
rect 11732 37996 11742 38052
rect 11442 37772 11452 37828
rect 11508 37772 15932 37828
rect 15988 37772 15998 37828
rect 26852 37772 27804 37828
rect 27860 37772 27870 37828
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 26852 37604 26908 37772
rect 22194 37548 22204 37604
rect 22260 37548 23996 37604
rect 24052 37548 26908 37604
rect 16146 37436 16156 37492
rect 16212 37436 17388 37492
rect 17444 37436 17454 37492
rect 27570 37436 27580 37492
rect 27636 37436 30268 37492
rect 30324 37436 31612 37492
rect 31668 37436 31678 37492
rect 31826 37436 31836 37492
rect 31892 37436 32396 37492
rect 32452 37436 34972 37492
rect 35028 37436 35038 37492
rect 25218 37324 25228 37380
rect 25284 37324 25788 37380
rect 25844 37324 28700 37380
rect 28756 37324 29484 37380
rect 29540 37324 30660 37380
rect 31378 37324 31388 37380
rect 31444 37324 32732 37380
rect 32788 37324 33740 37380
rect 33796 37324 33806 37380
rect 30604 37268 30660 37324
rect 19506 37212 19516 37268
rect 19572 37212 23548 37268
rect 23604 37212 25900 37268
rect 25956 37212 25966 37268
rect 27906 37212 27916 37268
rect 27972 37212 29820 37268
rect 29876 37212 29886 37268
rect 30604 37212 31500 37268
rect 31556 37212 33628 37268
rect 33684 37212 33694 37268
rect 11218 37100 11228 37156
rect 11284 37100 12908 37156
rect 12964 37100 12974 37156
rect 14802 36988 14812 37044
rect 14868 36988 15372 37044
rect 15428 36988 15708 37044
rect 15764 36988 15774 37044
rect 25330 36988 25340 37044
rect 25396 36988 27244 37044
rect 27300 36988 27310 37044
rect 15138 36876 15148 36932
rect 15204 36876 16156 36932
rect 16212 36876 16222 36932
rect 25890 36876 25900 36932
rect 25956 36876 29036 36932
rect 29092 36876 29820 36932
rect 29876 36876 31276 36932
rect 31332 36876 32508 36932
rect 32564 36876 32844 36932
rect 32900 36876 34076 36932
rect 34132 36876 34142 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 12562 36764 12572 36820
rect 12628 36764 13916 36820
rect 13972 36764 13982 36820
rect 23650 36764 23660 36820
rect 23716 36764 24668 36820
rect 24724 36764 26236 36820
rect 26292 36764 26302 36820
rect 12114 36652 12124 36708
rect 12180 36652 13468 36708
rect 13524 36652 13534 36708
rect 33170 36652 33180 36708
rect 33236 36652 35532 36708
rect 35588 36652 36540 36708
rect 36596 36652 36606 36708
rect 12898 36540 12908 36596
rect 12964 36540 13580 36596
rect 13636 36540 13646 36596
rect 26562 36540 26572 36596
rect 26628 36540 27580 36596
rect 27636 36540 27646 36596
rect 7522 36428 7532 36484
rect 7588 36428 9100 36484
rect 9156 36428 10780 36484
rect 10836 36428 11676 36484
rect 11732 36428 13132 36484
rect 13188 36428 15260 36484
rect 15316 36428 16492 36484
rect 16548 36428 16558 36484
rect 24210 36428 24220 36484
rect 24276 36428 25340 36484
rect 25396 36428 25406 36484
rect 29698 36428 29708 36484
rect 29764 36428 30716 36484
rect 30772 36428 30782 36484
rect 32050 36428 32060 36484
rect 32116 36428 33404 36484
rect 33460 36428 33470 36484
rect 0 36372 800 36400
rect 0 36316 4060 36372
rect 4116 36316 4126 36372
rect 18610 36316 18620 36372
rect 18676 36316 20524 36372
rect 20580 36316 21756 36372
rect 21812 36316 22988 36372
rect 23044 36316 23884 36372
rect 23940 36316 23950 36372
rect 26114 36316 26124 36372
rect 26180 36316 27692 36372
rect 27748 36316 27758 36372
rect 28466 36316 28476 36372
rect 28532 36316 29596 36372
rect 29652 36316 29662 36372
rect 30930 36316 30940 36372
rect 30996 36316 31948 36372
rect 32004 36316 32014 36372
rect 0 36288 800 36316
rect 26124 36260 26180 36316
rect 11890 36204 11900 36260
rect 11956 36204 12796 36260
rect 12852 36204 12862 36260
rect 15698 36204 15708 36260
rect 15764 36204 16716 36260
rect 16772 36204 16782 36260
rect 19618 36204 19628 36260
rect 19684 36204 20412 36260
rect 20468 36204 20478 36260
rect 20962 36204 20972 36260
rect 21028 36204 21532 36260
rect 21588 36204 26180 36260
rect 27692 36260 27748 36316
rect 27692 36204 29372 36260
rect 29428 36204 30268 36260
rect 30324 36204 30828 36260
rect 30884 36204 30894 36260
rect 34402 36204 34412 36260
rect 34468 36204 35756 36260
rect 35812 36204 35822 36260
rect 15922 36092 15932 36148
rect 15988 36092 16380 36148
rect 16436 36092 18060 36148
rect 18116 36092 18126 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 13906 35980 13916 36036
rect 13972 35980 18620 36036
rect 18676 35980 18686 36036
rect 20402 35980 20412 36036
rect 20468 35980 21532 36036
rect 21588 35980 22092 36036
rect 22148 35980 22158 36036
rect 9538 35868 9548 35924
rect 9604 35868 11340 35924
rect 11396 35868 11406 35924
rect 18274 35868 18284 35924
rect 18340 35868 19180 35924
rect 19236 35868 19246 35924
rect 27346 35868 27356 35924
rect 27412 35868 28364 35924
rect 28420 35868 28430 35924
rect 15698 35756 15708 35812
rect 15764 35756 19628 35812
rect 19684 35756 19694 35812
rect 10994 35644 11004 35700
rect 11060 35644 11452 35700
rect 11508 35644 16492 35700
rect 16548 35644 16828 35700
rect 16884 35644 16894 35700
rect 17826 35644 17836 35700
rect 17892 35644 18284 35700
rect 18340 35644 19740 35700
rect 19796 35644 19806 35700
rect 20290 35644 20300 35700
rect 20356 35644 21308 35700
rect 21364 35644 21374 35700
rect 21746 35644 21756 35700
rect 21812 35644 24220 35700
rect 24276 35644 24286 35700
rect 26674 35644 26684 35700
rect 26740 35644 27972 35700
rect 30818 35644 30828 35700
rect 30884 35644 32060 35700
rect 32116 35644 33740 35700
rect 33796 35644 33806 35700
rect 27916 35588 27972 35644
rect 13906 35532 13916 35588
rect 13972 35532 14476 35588
rect 14532 35532 17388 35588
rect 17444 35532 17454 35588
rect 17612 35532 17948 35588
rect 18004 35532 18014 35588
rect 20738 35532 20748 35588
rect 20804 35532 22316 35588
rect 22372 35532 25788 35588
rect 25844 35532 25854 35588
rect 27906 35532 27916 35588
rect 27972 35532 28812 35588
rect 28868 35532 30268 35588
rect 30324 35532 30492 35588
rect 30548 35532 33628 35588
rect 33684 35532 34300 35588
rect 34356 35532 34366 35588
rect 17612 35476 17668 35532
rect 15026 35420 15036 35476
rect 15092 35420 15260 35476
rect 15316 35420 15708 35476
rect 15764 35420 15774 35476
rect 17154 35420 17164 35476
rect 17220 35420 17668 35476
rect 33282 35420 33292 35476
rect 33348 35420 33852 35476
rect 33908 35420 34860 35476
rect 34916 35420 34926 35476
rect 11676 35308 12236 35364
rect 12292 35308 12302 35364
rect 16482 35308 16492 35364
rect 16548 35308 19852 35364
rect 19908 35308 20972 35364
rect 21028 35308 21038 35364
rect 21298 35308 21308 35364
rect 21364 35308 24388 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 11676 35252 11732 35308
rect 24332 35252 24388 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 11666 35196 11676 35252
rect 11732 35196 11742 35252
rect 16034 35196 16044 35252
rect 16100 35196 16380 35252
rect 16436 35196 16446 35252
rect 24322 35196 24332 35252
rect 24388 35196 24398 35252
rect 14914 35084 14924 35140
rect 14980 35084 15260 35140
rect 15316 35084 15326 35140
rect 16156 35084 18396 35140
rect 18452 35084 19180 35140
rect 19236 35084 19246 35140
rect 20738 35084 20748 35140
rect 20804 35084 22652 35140
rect 22708 35084 22718 35140
rect 16156 35028 16212 35084
rect 12450 34972 12460 35028
rect 12516 34972 16212 35028
rect 16370 34972 16380 35028
rect 16436 34972 18844 35028
rect 18900 34972 18910 35028
rect 20626 34972 20636 35028
rect 20692 34972 21980 35028
rect 22036 34972 22428 35028
rect 22484 34972 22988 35028
rect 23044 34972 23054 35028
rect 24546 34972 24556 35028
rect 24612 34972 25228 35028
rect 25284 34972 25294 35028
rect 14018 34860 14028 34916
rect 14084 34860 14476 34916
rect 14532 34860 14542 34916
rect 14690 34860 14700 34916
rect 14756 34860 16044 34916
rect 16100 34860 16110 34916
rect 16482 34860 16492 34916
rect 16548 34860 16828 34916
rect 16884 34860 16894 34916
rect 17490 34860 17500 34916
rect 17556 34860 18172 34916
rect 18228 34860 18732 34916
rect 18788 34860 18798 34916
rect 20962 34860 20972 34916
rect 21028 34860 21756 34916
rect 21812 34860 23436 34916
rect 23492 34860 23502 34916
rect 24210 34860 24220 34916
rect 24276 34860 25676 34916
rect 25732 34860 29820 34916
rect 29876 34860 29886 34916
rect 30818 34860 30828 34916
rect 30884 34860 31388 34916
rect 31444 34860 33964 34916
rect 34020 34860 34030 34916
rect 14802 34748 14812 34804
rect 14868 34748 15820 34804
rect 15876 34748 15886 34804
rect 16258 34748 16268 34804
rect 16324 34748 20300 34804
rect 20356 34748 20366 34804
rect 24546 34748 24556 34804
rect 24612 34748 25228 34804
rect 25284 34748 26572 34804
rect 26628 34748 26638 34804
rect 26572 34692 26628 34748
rect 9090 34636 9100 34692
rect 9156 34636 10108 34692
rect 10164 34636 10174 34692
rect 13010 34636 13020 34692
rect 13076 34636 13692 34692
rect 13748 34636 14700 34692
rect 14756 34636 14766 34692
rect 15250 34636 15260 34692
rect 15316 34636 16380 34692
rect 16436 34636 16446 34692
rect 18610 34636 18620 34692
rect 18676 34636 18686 34692
rect 26572 34636 26908 34692
rect 26964 34636 26974 34692
rect 27346 34636 27356 34692
rect 27412 34636 28364 34692
rect 28420 34636 29372 34692
rect 29428 34636 30940 34692
rect 30996 34636 31836 34692
rect 31892 34636 31902 34692
rect 18620 34580 18676 34636
rect 14466 34524 14476 34580
rect 14532 34524 18676 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 26852 34468 26908 34636
rect 14690 34412 14700 34468
rect 14756 34412 15596 34468
rect 15652 34412 15662 34468
rect 22418 34412 22428 34468
rect 22484 34412 23436 34468
rect 23492 34412 24780 34468
rect 24836 34412 24846 34468
rect 26852 34412 29428 34468
rect 29372 34356 29428 34412
rect 7410 34300 7420 34356
rect 7476 34300 8540 34356
rect 8596 34300 8606 34356
rect 16930 34300 16940 34356
rect 16996 34300 17724 34356
rect 17780 34300 18508 34356
rect 18564 34300 18574 34356
rect 23314 34300 23324 34356
rect 23380 34300 23660 34356
rect 23716 34300 25116 34356
rect 25172 34300 25182 34356
rect 27234 34300 27244 34356
rect 27300 34300 27916 34356
rect 27972 34300 27982 34356
rect 29362 34300 29372 34356
rect 29428 34300 30828 34356
rect 30884 34300 30894 34356
rect 15698 34188 15708 34244
rect 15764 34188 17388 34244
rect 17444 34188 18844 34244
rect 18900 34188 19180 34244
rect 19236 34188 19246 34244
rect 22754 34188 22764 34244
rect 22820 34188 25676 34244
rect 25732 34188 25742 34244
rect 26852 34188 28028 34244
rect 28084 34188 28094 34244
rect 24668 34132 24724 34188
rect 26852 34132 26908 34188
rect 8082 34076 8092 34132
rect 8148 34076 8876 34132
rect 8932 34076 8942 34132
rect 9202 34076 9212 34132
rect 9268 34076 10108 34132
rect 10164 34076 10174 34132
rect 11890 34076 11900 34132
rect 11956 34076 12684 34132
rect 12740 34076 12750 34132
rect 13906 34076 13916 34132
rect 13972 34076 15036 34132
rect 15092 34076 15596 34132
rect 15652 34076 15662 34132
rect 22306 34076 22316 34132
rect 22372 34076 22652 34132
rect 22708 34076 24108 34132
rect 24164 34076 24174 34132
rect 24658 34076 24668 34132
rect 24724 34076 24734 34132
rect 24882 34076 24892 34132
rect 24948 34076 25228 34132
rect 25284 34076 25294 34132
rect 26226 34076 26236 34132
rect 26292 34076 26908 34132
rect 27122 34076 27132 34132
rect 27188 34076 28140 34132
rect 28196 34076 28206 34132
rect 29810 34076 29820 34132
rect 29876 34076 30492 34132
rect 30548 34076 30558 34132
rect 33618 34076 33628 34132
rect 33684 34076 35084 34132
rect 35140 34076 35150 34132
rect 10322 33964 10332 34020
rect 10388 33964 11452 34020
rect 11508 33964 11518 34020
rect 12002 33964 12012 34020
rect 12068 33964 12796 34020
rect 12852 33964 12862 34020
rect 15092 33964 16604 34020
rect 16660 33964 16670 34020
rect 22082 33964 22092 34020
rect 22148 33964 24332 34020
rect 24388 33964 24398 34020
rect 26114 33964 26124 34020
rect 26180 33964 26190 34020
rect 26450 33964 26460 34020
rect 26516 33964 27412 34020
rect 11452 33908 11508 33964
rect 15092 33908 15148 33964
rect 3938 33852 3948 33908
rect 4004 33852 6468 33908
rect 11452 33852 15148 33908
rect 23986 33852 23996 33908
rect 24052 33852 24062 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 6412 33684 6468 33852
rect 14018 33740 14028 33796
rect 14084 33740 14588 33796
rect 14644 33740 14654 33796
rect 23996 33684 24052 33852
rect 26124 33796 26180 33964
rect 26796 33852 27132 33908
rect 27188 33852 27198 33908
rect 26796 33796 26852 33852
rect 27356 33796 27412 33964
rect 32050 33852 32060 33908
rect 32116 33852 32508 33908
rect 32564 33852 32574 33908
rect 26124 33740 26852 33796
rect 27346 33740 27356 33796
rect 27412 33740 27916 33796
rect 27972 33740 27982 33796
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 6402 33628 6412 33684
rect 6468 33628 7532 33684
rect 7588 33628 7598 33684
rect 23996 33628 26460 33684
rect 26516 33628 26526 33684
rect 30370 33628 30380 33684
rect 30436 33628 32396 33684
rect 32452 33628 33740 33684
rect 33796 33628 33806 33684
rect 6626 33516 6636 33572
rect 6692 33516 6972 33572
rect 7028 33516 7038 33572
rect 9762 33516 9772 33572
rect 9828 33516 10556 33572
rect 10612 33516 10622 33572
rect 13682 33516 13692 33572
rect 13748 33516 15148 33572
rect 16594 33516 16604 33572
rect 16660 33516 17836 33572
rect 17892 33516 17902 33572
rect 4274 33404 4284 33460
rect 4340 33404 6188 33460
rect 6244 33404 6254 33460
rect 15092 33348 15148 33516
rect 17042 33404 17052 33460
rect 17108 33404 19068 33460
rect 19124 33404 19134 33460
rect 23996 33348 24052 33628
rect 26114 33516 26124 33572
rect 26180 33516 27804 33572
rect 27860 33516 27870 33572
rect 32722 33516 32732 33572
rect 32788 33516 33068 33572
rect 33124 33516 33134 33572
rect 32498 33404 32508 33460
rect 32564 33404 33628 33460
rect 33684 33404 33694 33460
rect 7858 33292 7868 33348
rect 7924 33292 8876 33348
rect 8932 33292 10108 33348
rect 10164 33292 10174 33348
rect 13794 33292 13804 33348
rect 13860 33292 14700 33348
rect 14756 33292 14766 33348
rect 15092 33292 16604 33348
rect 16660 33292 16670 33348
rect 23986 33292 23996 33348
rect 24052 33292 24062 33348
rect 31490 33292 31500 33348
rect 31556 33292 32172 33348
rect 32228 33292 32788 33348
rect 32946 33292 32956 33348
rect 33012 33292 35084 33348
rect 35140 33292 35150 33348
rect 32732 33236 32788 33292
rect 13682 33180 13692 33236
rect 13748 33180 16716 33236
rect 16772 33180 18396 33236
rect 18452 33180 18462 33236
rect 21858 33180 21868 33236
rect 21924 33180 24220 33236
rect 24276 33180 24286 33236
rect 30482 33180 30492 33236
rect 30548 33180 32284 33236
rect 32340 33180 32350 33236
rect 32732 33180 33628 33236
rect 33684 33180 34972 33236
rect 35028 33180 35038 33236
rect 6066 33068 6076 33124
rect 6132 33068 8652 33124
rect 8708 33068 8718 33124
rect 10098 33068 10108 33124
rect 10164 33068 11116 33124
rect 11172 33068 11676 33124
rect 11732 33068 11742 33124
rect 18834 33068 18844 33124
rect 18900 33068 19180 33124
rect 19236 33068 19246 33124
rect 19394 33068 19404 33124
rect 19460 33068 19964 33124
rect 20020 33068 21980 33124
rect 22036 33068 22046 33124
rect 26226 33068 26236 33124
rect 26292 33068 27356 33124
rect 27412 33068 27422 33124
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 9090 32732 9100 32788
rect 9156 32732 9884 32788
rect 9940 32732 9950 32788
rect 12562 32732 12572 32788
rect 12628 32732 13580 32788
rect 13636 32732 13646 32788
rect 30818 32732 30828 32788
rect 30884 32732 32732 32788
rect 32788 32732 34188 32788
rect 34244 32732 34254 32788
rect 8978 32620 8988 32676
rect 9044 32620 10108 32676
rect 10164 32620 10174 32676
rect 10882 32620 10892 32676
rect 10948 32620 11452 32676
rect 11508 32620 11518 32676
rect 12786 32620 12796 32676
rect 12852 32620 13692 32676
rect 13748 32620 13758 32676
rect 18386 32620 18396 32676
rect 18452 32620 19292 32676
rect 19348 32620 19358 32676
rect 24098 32620 24108 32676
rect 24164 32620 26908 32676
rect 26964 32620 26974 32676
rect 28018 32620 28028 32676
rect 28084 32620 28476 32676
rect 28532 32620 28542 32676
rect 33394 32620 33404 32676
rect 33460 32620 34076 32676
rect 34132 32620 34142 32676
rect 9874 32508 9884 32564
rect 9940 32508 11116 32564
rect 11172 32508 11182 32564
rect 17826 32508 17836 32564
rect 17892 32508 19404 32564
rect 19460 32508 19470 32564
rect 33170 32508 33180 32564
rect 33236 32508 33628 32564
rect 33684 32508 34188 32564
rect 34244 32508 34254 32564
rect 6066 32396 6076 32452
rect 6132 32396 7196 32452
rect 7252 32396 7262 32452
rect 20178 32396 20188 32452
rect 20244 32396 20972 32452
rect 21028 32396 21038 32452
rect 21858 32396 21868 32452
rect 21924 32396 22204 32452
rect 22260 32396 22270 32452
rect 27346 32396 27356 32452
rect 27412 32396 28140 32452
rect 28196 32396 28206 32452
rect 22418 32172 22428 32228
rect 22484 32172 22764 32228
rect 22820 32172 24108 32228
rect 24164 32172 24174 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 5954 32060 5964 32116
rect 6020 32060 6300 32116
rect 6356 32060 6860 32116
rect 6916 32060 6926 32116
rect 12562 32060 12572 32116
rect 12628 32060 13468 32116
rect 13524 32060 14140 32116
rect 14196 32060 14206 32116
rect 30930 32060 30940 32116
rect 30996 32060 31500 32116
rect 31556 32060 31566 32116
rect 21970 31948 21980 32004
rect 22036 31948 22652 32004
rect 22708 31948 22718 32004
rect 31714 31948 31724 32004
rect 31780 31948 32508 32004
rect 32564 31948 33180 32004
rect 33236 31948 33246 32004
rect 8194 31836 8204 31892
rect 8260 31836 9884 31892
rect 9940 31836 9950 31892
rect 13906 31836 13916 31892
rect 13972 31836 14924 31892
rect 14980 31836 14990 31892
rect 24658 31836 24668 31892
rect 24724 31836 26348 31892
rect 26404 31836 26414 31892
rect 27010 31836 27020 31892
rect 27076 31836 27692 31892
rect 27748 31836 27758 31892
rect 28018 31836 28028 31892
rect 28084 31836 30492 31892
rect 30548 31836 30558 31892
rect 30930 31836 30940 31892
rect 30996 31836 31388 31892
rect 31444 31836 32060 31892
rect 32116 31836 32126 31892
rect 30492 31780 30548 31836
rect 9538 31724 9548 31780
rect 9604 31724 13300 31780
rect 14690 31724 14700 31780
rect 14756 31724 17276 31780
rect 17332 31724 17342 31780
rect 19506 31724 19516 31780
rect 19572 31724 20524 31780
rect 20580 31724 20590 31780
rect 20738 31724 20748 31780
rect 20804 31724 22428 31780
rect 22484 31724 23436 31780
rect 23492 31724 23502 31780
rect 24434 31724 24444 31780
rect 24500 31724 25676 31780
rect 25732 31724 26572 31780
rect 26628 31724 26638 31780
rect 26786 31724 26796 31780
rect 26852 31724 27804 31780
rect 27860 31724 27870 31780
rect 28242 31724 28252 31780
rect 28308 31724 29148 31780
rect 29204 31724 29214 31780
rect 30492 31724 31836 31780
rect 31892 31724 31902 31780
rect 13244 31668 13300 31724
rect 41200 31668 42000 31696
rect 2034 31612 2044 31668
rect 2100 31612 7308 31668
rect 7364 31612 7756 31668
rect 7812 31612 7822 31668
rect 8866 31612 8876 31668
rect 8932 31612 10108 31668
rect 10164 31612 10174 31668
rect 11554 31612 11564 31668
rect 11620 31612 12124 31668
rect 12180 31612 13020 31668
rect 13076 31612 13086 31668
rect 13244 31612 13468 31668
rect 13524 31612 13916 31668
rect 13972 31612 13982 31668
rect 14354 31612 14364 31668
rect 14420 31612 15596 31668
rect 15652 31612 15662 31668
rect 16818 31612 16828 31668
rect 16884 31612 18396 31668
rect 18452 31612 19292 31668
rect 19348 31612 19740 31668
rect 19796 31612 19806 31668
rect 22194 31612 22204 31668
rect 22260 31612 23212 31668
rect 23268 31612 23278 31668
rect 26002 31612 26012 31668
rect 26068 31612 26078 31668
rect 26898 31612 26908 31668
rect 26964 31612 27580 31668
rect 27636 31612 27646 31668
rect 28578 31612 28588 31668
rect 28644 31612 29260 31668
rect 29316 31612 29326 31668
rect 29810 31612 29820 31668
rect 29876 31612 30604 31668
rect 30660 31612 31612 31668
rect 31668 31612 31678 31668
rect 39554 31612 39564 31668
rect 39620 31612 40012 31668
rect 40068 31612 42000 31668
rect 26012 31556 26068 31612
rect 41200 31584 42000 31612
rect 1698 31500 1708 31556
rect 1764 31500 2492 31556
rect 2548 31500 2558 31556
rect 3266 31500 3276 31556
rect 3332 31500 5740 31556
rect 5796 31500 5806 31556
rect 18722 31500 18732 31556
rect 18788 31500 19516 31556
rect 19572 31500 19582 31556
rect 23314 31500 23324 31556
rect 23380 31500 23390 31556
rect 26012 31500 27244 31556
rect 27300 31500 27310 31556
rect 33058 31500 33068 31556
rect 33124 31500 34076 31556
rect 34132 31500 34142 31556
rect 23324 31444 23380 31500
rect 23324 31388 30716 31444
rect 30772 31388 31164 31444
rect 31220 31388 31230 31444
rect 31490 31388 31500 31444
rect 31556 31388 33516 31444
rect 33572 31388 39900 31444
rect 39956 31388 39966 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 8754 31276 8764 31332
rect 8820 31276 9548 31332
rect 9604 31276 9614 31332
rect 13682 31164 13692 31220
rect 13748 31164 14924 31220
rect 14980 31164 15372 31220
rect 15428 31164 15438 31220
rect 16706 31164 16716 31220
rect 16772 31164 18284 31220
rect 18340 31164 18350 31220
rect 19506 31164 19516 31220
rect 19572 31164 20636 31220
rect 20692 31164 20702 31220
rect 26114 31164 26124 31220
rect 26180 31164 26796 31220
rect 26852 31164 26862 31220
rect 31602 31164 31612 31220
rect 31668 31164 32844 31220
rect 32900 31164 32910 31220
rect 2818 31052 2828 31108
rect 2884 31052 6524 31108
rect 6580 31052 6590 31108
rect 7410 31052 7420 31108
rect 7476 31052 8540 31108
rect 8596 31052 9212 31108
rect 9268 31052 9660 31108
rect 9716 31052 9726 31108
rect 13458 31052 13468 31108
rect 13524 31052 14028 31108
rect 14084 31052 14094 31108
rect 14802 31052 14812 31108
rect 14868 31052 18508 31108
rect 18564 31052 18574 31108
rect 32162 31052 32172 31108
rect 32228 31052 33292 31108
rect 33348 31052 33358 31108
rect 0 30996 800 31024
rect 6524 30996 6580 31052
rect 41200 30996 42000 31024
rect 0 30940 1708 30996
rect 1764 30940 1774 30996
rect 6524 30940 7980 30996
rect 8036 30940 8652 30996
rect 8708 30940 9324 30996
rect 9380 30940 9390 30996
rect 11442 30940 11452 30996
rect 11508 30940 12124 30996
rect 12180 30940 12190 30996
rect 15474 30940 15484 30996
rect 15540 30940 17500 30996
rect 17556 30940 17566 30996
rect 18162 30940 18172 30996
rect 18228 30940 18956 30996
rect 19012 30940 19022 30996
rect 26002 30940 26012 30996
rect 26068 30940 26684 30996
rect 26740 30940 26750 30996
rect 32386 30940 32396 30996
rect 32452 30940 33740 30996
rect 33796 30940 34860 30996
rect 34916 30940 34926 30996
rect 40226 30940 40236 30996
rect 40292 30940 42000 30996
rect 0 30912 800 30940
rect 41200 30912 42000 30940
rect 12786 30828 12796 30884
rect 12852 30828 15260 30884
rect 15316 30828 15326 30884
rect 16594 30828 16604 30884
rect 16660 30828 17164 30884
rect 17220 30828 17230 30884
rect 18050 30828 18060 30884
rect 18116 30828 18732 30884
rect 18788 30828 18798 30884
rect 27458 30828 27468 30884
rect 27524 30828 29260 30884
rect 29316 30828 29326 30884
rect 32050 30828 32060 30884
rect 32116 30828 33068 30884
rect 33124 30828 33134 30884
rect 11778 30716 11788 30772
rect 11844 30716 12460 30772
rect 12516 30716 12526 30772
rect 30594 30716 30604 30772
rect 30660 30716 31948 30772
rect 32004 30716 32014 30772
rect 11218 30604 11228 30660
rect 11284 30604 22316 30660
rect 22372 30604 23324 30660
rect 23380 30604 23390 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 11228 30436 11284 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 8316 30380 11284 30436
rect 14242 30380 14252 30436
rect 14308 30380 18620 30436
rect 18676 30380 18686 30436
rect 19170 30380 19180 30436
rect 19236 30380 21308 30436
rect 21364 30380 21374 30436
rect 32274 30380 32284 30436
rect 32340 30380 35420 30436
rect 35476 30380 35486 30436
rect 0 30324 800 30352
rect 8316 30324 8372 30380
rect 0 30268 2212 30324
rect 0 30240 800 30268
rect 2156 30212 2212 30268
rect 8092 30268 8372 30324
rect 9762 30268 9772 30324
rect 9828 30268 11452 30324
rect 11508 30268 11518 30324
rect 17378 30268 17388 30324
rect 17444 30268 18508 30324
rect 18564 30268 18574 30324
rect 33394 30268 33404 30324
rect 33460 30268 35644 30324
rect 35700 30268 39228 30324
rect 39284 30268 39294 30324
rect 8092 30212 8148 30268
rect 2146 30156 2156 30212
rect 2212 30156 2222 30212
rect 6066 30156 6076 30212
rect 6132 30156 6748 30212
rect 6804 30156 8148 30212
rect 8306 30156 8316 30212
rect 8372 30156 10220 30212
rect 10276 30156 10286 30212
rect 10434 30156 10444 30212
rect 10500 30156 11004 30212
rect 11060 30156 11900 30212
rect 11956 30156 11966 30212
rect 12226 30156 12236 30212
rect 12292 30156 14028 30212
rect 14084 30156 14094 30212
rect 14466 30156 14476 30212
rect 14532 30156 15484 30212
rect 15540 30156 15550 30212
rect 17154 30156 17164 30212
rect 17220 30156 18284 30212
rect 18340 30156 18350 30212
rect 18722 30156 18732 30212
rect 18788 30156 20076 30212
rect 20132 30156 22092 30212
rect 22148 30156 22158 30212
rect 25890 30156 25900 30212
rect 25956 30156 27916 30212
rect 27972 30156 29148 30212
rect 29204 30156 29214 30212
rect 31266 30156 31276 30212
rect 31332 30156 32396 30212
rect 32452 30156 33180 30212
rect 33236 30156 33246 30212
rect 6514 30044 6524 30100
rect 6580 30044 7308 30100
rect 7364 30044 7374 30100
rect 16146 30044 16156 30100
rect 16212 30044 16940 30100
rect 16996 30044 17006 30100
rect 17714 30044 17724 30100
rect 17780 30044 18172 30100
rect 18228 30044 18238 30100
rect 19180 30044 22204 30100
rect 22260 30044 22270 30100
rect 24546 30044 24556 30100
rect 24612 30044 25004 30100
rect 25060 30044 26348 30100
rect 26404 30044 26572 30100
rect 26628 30044 26638 30100
rect 26898 30044 26908 30100
rect 26964 30044 27804 30100
rect 27860 30044 27870 30100
rect 32498 30044 32508 30100
rect 32564 30044 34524 30100
rect 34580 30044 34590 30100
rect 19180 29988 19236 30044
rect 5170 29932 5180 29988
rect 5236 29932 6300 29988
rect 6356 29932 8540 29988
rect 8596 29932 9548 29988
rect 9604 29932 9614 29988
rect 14578 29932 14588 29988
rect 14644 29932 19236 29988
rect 19394 29932 19404 29988
rect 19460 29932 20300 29988
rect 20356 29932 20366 29988
rect 20514 29932 20524 29988
rect 20580 29932 20972 29988
rect 21028 29932 24220 29988
rect 24276 29932 24286 29988
rect 24658 29932 24668 29988
rect 24724 29932 25788 29988
rect 25844 29932 25854 29988
rect 14130 29820 14140 29876
rect 14196 29820 17052 29876
rect 17108 29820 17118 29876
rect 17388 29820 17612 29876
rect 17668 29820 17678 29876
rect 22082 29820 22092 29876
rect 22148 29820 29596 29876
rect 29652 29820 29662 29876
rect 8082 29708 8092 29764
rect 8148 29708 10220 29764
rect 10276 29708 10286 29764
rect 9314 29596 9324 29652
rect 9380 29596 10444 29652
rect 10500 29596 10510 29652
rect 16370 29596 16380 29652
rect 16436 29596 17164 29652
rect 17220 29596 17230 29652
rect 6626 29484 6636 29540
rect 6692 29484 6702 29540
rect 7634 29484 7644 29540
rect 7700 29484 8876 29540
rect 8932 29484 8942 29540
rect 6636 29428 6692 29484
rect 17388 29428 17444 29820
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 19506 29708 19516 29764
rect 19572 29708 19582 29764
rect 24210 29708 24220 29764
rect 24276 29708 26012 29764
rect 26068 29708 26078 29764
rect 19516 29652 19572 29708
rect 17938 29596 17948 29652
rect 18004 29596 18014 29652
rect 19282 29596 19292 29652
rect 19348 29596 20412 29652
rect 20468 29596 21644 29652
rect 21700 29596 22540 29652
rect 22596 29596 22606 29652
rect 26852 29596 30828 29652
rect 30884 29596 32060 29652
rect 32116 29596 34412 29652
rect 34468 29596 37100 29652
rect 37156 29596 37166 29652
rect 17948 29428 18004 29596
rect 19058 29484 19068 29540
rect 19124 29484 20188 29540
rect 20244 29484 20254 29540
rect 5618 29372 5628 29428
rect 5684 29372 6692 29428
rect 10098 29372 10108 29428
rect 10164 29372 10556 29428
rect 10612 29372 10622 29428
rect 16146 29372 16156 29428
rect 16212 29372 16828 29428
rect 16884 29372 16894 29428
rect 17378 29372 17388 29428
rect 17444 29372 17454 29428
rect 17602 29372 17612 29428
rect 17668 29372 18004 29428
rect 19954 29372 19964 29428
rect 20020 29372 20300 29428
rect 20356 29372 20366 29428
rect 25554 29372 25564 29428
rect 25620 29372 26348 29428
rect 26404 29372 26414 29428
rect 26852 29316 26908 29596
rect 28578 29484 28588 29540
rect 28644 29484 31388 29540
rect 31444 29484 32508 29540
rect 32564 29484 32574 29540
rect 33954 29372 33964 29428
rect 34020 29372 35196 29428
rect 35252 29372 35262 29428
rect 37426 29372 37436 29428
rect 37492 29372 39004 29428
rect 39060 29372 39070 29428
rect 6066 29260 6076 29316
rect 6132 29260 6636 29316
rect 6692 29260 6702 29316
rect 15092 29260 16268 29316
rect 16324 29260 20972 29316
rect 21028 29260 21038 29316
rect 25218 29260 25228 29316
rect 25284 29260 25788 29316
rect 25844 29260 26908 29316
rect 30370 29260 30380 29316
rect 30436 29260 31724 29316
rect 31780 29260 34972 29316
rect 35028 29260 35868 29316
rect 35924 29260 35934 29316
rect 0 28980 800 29008
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 15092 28980 15148 29260
rect 25330 29148 25340 29204
rect 25396 29148 25900 29204
rect 25956 29148 25966 29204
rect 32722 29148 32732 29204
rect 32788 29148 33516 29204
rect 33572 29148 39900 29204
rect 39956 29148 39966 29204
rect 32498 29036 32508 29092
rect 32564 29036 34748 29092
rect 34804 29036 34814 29092
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 41200 28980 42000 29008
rect 0 28924 1708 28980
rect 1764 28924 2492 28980
rect 2548 28924 2558 28980
rect 10210 28924 10220 28980
rect 10276 28924 11900 28980
rect 11956 28924 15148 28980
rect 32946 28924 32956 28980
rect 33012 28924 33292 28980
rect 33348 28924 35028 28980
rect 40114 28924 40124 28980
rect 40180 28924 42000 28980
rect 0 28896 800 28924
rect 34972 28868 35028 28924
rect 41200 28896 42000 28924
rect 2034 28812 2044 28868
rect 2100 28812 8652 28868
rect 8708 28812 8718 28868
rect 9874 28812 9884 28868
rect 9940 28812 10556 28868
rect 10612 28812 11340 28868
rect 11396 28812 14140 28868
rect 14196 28812 14206 28868
rect 16706 28812 16716 28868
rect 16772 28812 17724 28868
rect 17780 28812 17790 28868
rect 34972 28812 35532 28868
rect 35588 28812 35598 28868
rect 2930 28700 2940 28756
rect 2996 28700 6860 28756
rect 6916 28700 7308 28756
rect 7364 28700 7644 28756
rect 7700 28700 7710 28756
rect 8306 28700 8316 28756
rect 8372 28700 9772 28756
rect 9828 28700 10108 28756
rect 10164 28700 11004 28756
rect 11060 28700 11070 28756
rect 15474 28700 15484 28756
rect 15540 28700 16828 28756
rect 16884 28700 17948 28756
rect 18004 28700 18014 28756
rect 18610 28700 18620 28756
rect 18676 28700 19964 28756
rect 20020 28700 20030 28756
rect 26852 28700 27356 28756
rect 27412 28700 30716 28756
rect 30772 28700 31500 28756
rect 31556 28700 31566 28756
rect 33170 28700 33180 28756
rect 33236 28700 33964 28756
rect 34020 28700 35420 28756
rect 35476 28700 37436 28756
rect 37492 28700 37502 28756
rect 8194 28588 8204 28644
rect 8260 28588 8764 28644
rect 8820 28588 8830 28644
rect 10546 28588 10556 28644
rect 10612 28588 11452 28644
rect 11508 28588 12460 28644
rect 12516 28588 12526 28644
rect 14354 28588 14364 28644
rect 14420 28588 15148 28644
rect 15204 28588 15214 28644
rect 16258 28476 16268 28532
rect 16324 28476 17276 28532
rect 17332 28476 17342 28532
rect 2146 28364 2156 28420
rect 2212 28364 2222 28420
rect 4274 28364 4284 28420
rect 4340 28364 5964 28420
rect 6020 28364 6030 28420
rect 10770 28364 10780 28420
rect 10836 28364 17164 28420
rect 17220 28364 18396 28420
rect 18452 28364 18462 28420
rect 19170 28364 19180 28420
rect 19236 28364 19628 28420
rect 19684 28364 19694 28420
rect 0 28308 800 28336
rect 2156 28308 2212 28364
rect 26852 28308 26908 28700
rect 29138 28588 29148 28644
rect 29204 28588 29820 28644
rect 29876 28588 30380 28644
rect 30436 28588 32004 28644
rect 32162 28588 32172 28644
rect 32228 28588 33068 28644
rect 33124 28588 33134 28644
rect 34290 28588 34300 28644
rect 34356 28588 36316 28644
rect 36372 28588 36382 28644
rect 37090 28588 37100 28644
rect 37156 28588 37548 28644
rect 37604 28588 37614 28644
rect 31948 28532 32004 28588
rect 27010 28476 27020 28532
rect 27076 28476 27804 28532
rect 27860 28476 31052 28532
rect 31108 28476 31724 28532
rect 31780 28476 31790 28532
rect 31948 28476 32508 28532
rect 32564 28476 32574 28532
rect 33394 28476 33404 28532
rect 33460 28476 34636 28532
rect 34692 28476 34702 28532
rect 34402 28364 34412 28420
rect 34468 28364 36092 28420
rect 36148 28364 36158 28420
rect 41200 28308 42000 28336
rect 0 28252 2212 28308
rect 26338 28252 26348 28308
rect 26404 28252 26908 28308
rect 39666 28252 39676 28308
rect 39732 28252 40236 28308
rect 40292 28252 42000 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 41200 28224 42000 28252
rect 5842 28140 5852 28196
rect 5908 28140 10444 28196
rect 10500 28140 10510 28196
rect 6738 28028 6748 28084
rect 6804 28028 7532 28084
rect 7588 28028 7598 28084
rect 9650 28028 9660 28084
rect 9716 28028 10332 28084
rect 10388 28028 10398 28084
rect 15922 28028 15932 28084
rect 15988 28028 16604 28084
rect 16660 28028 18284 28084
rect 18340 28028 18350 28084
rect 23762 28028 23772 28084
rect 23828 28028 25116 28084
rect 25172 28028 25182 28084
rect 29698 28028 29708 28084
rect 29764 28028 30716 28084
rect 30772 28028 30782 28084
rect 30930 28028 30940 28084
rect 30996 28028 32396 28084
rect 32452 28028 32956 28084
rect 33012 28028 33022 28084
rect 3826 27804 3836 27860
rect 3892 27804 6188 27860
rect 6244 27804 7084 27860
rect 7140 27804 7150 27860
rect 19058 27804 19068 27860
rect 19124 27804 21196 27860
rect 21252 27804 22652 27860
rect 22708 27804 24780 27860
rect 24836 27804 26572 27860
rect 26628 27804 27580 27860
rect 27636 27804 28588 27860
rect 28644 27804 28654 27860
rect 29586 27804 29596 27860
rect 29652 27804 30380 27860
rect 30436 27804 31164 27860
rect 31220 27804 31948 27860
rect 32004 27804 32014 27860
rect 32610 27804 32620 27860
rect 32676 27804 33180 27860
rect 33236 27804 33740 27860
rect 33796 27804 33806 27860
rect 12898 27692 12908 27748
rect 12964 27692 13356 27748
rect 13412 27692 15932 27748
rect 15988 27692 15998 27748
rect 22978 27692 22988 27748
rect 23044 27692 25340 27748
rect 25396 27692 26684 27748
rect 26740 27692 26750 27748
rect 30594 27692 30604 27748
rect 30660 27692 31500 27748
rect 31556 27692 32172 27748
rect 32228 27692 32238 27748
rect 8082 27580 8092 27636
rect 8148 27580 14812 27636
rect 14868 27580 14878 27636
rect 21970 27580 21980 27636
rect 22036 27580 22876 27636
rect 22932 27580 22942 27636
rect 32274 27580 32284 27636
rect 32340 27580 32732 27636
rect 32788 27580 32798 27636
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 26674 27356 26684 27412
rect 26740 27356 28700 27412
rect 28756 27356 28766 27412
rect 9202 27244 9212 27300
rect 9268 27244 9884 27300
rect 9940 27244 10444 27300
rect 10500 27244 10510 27300
rect 29820 27244 33516 27300
rect 33572 27244 34748 27300
rect 34804 27244 34814 27300
rect 29820 27188 29876 27244
rect 8530 27132 8540 27188
rect 8596 27132 18396 27188
rect 18452 27132 18732 27188
rect 18788 27132 18798 27188
rect 24770 27132 24780 27188
rect 24836 27132 25452 27188
rect 25508 27132 25518 27188
rect 27458 27132 27468 27188
rect 27524 27132 29820 27188
rect 29876 27132 29886 27188
rect 31938 27132 31948 27188
rect 32004 27132 33404 27188
rect 33460 27132 33470 27188
rect 19058 27020 19068 27076
rect 19124 27020 19404 27076
rect 19460 27020 25900 27076
rect 25956 27020 26236 27076
rect 26292 27020 29484 27076
rect 29540 27020 29550 27076
rect 6290 26908 6300 26964
rect 6356 26908 11452 26964
rect 11508 26908 12348 26964
rect 12404 26908 16940 26964
rect 16996 26908 17388 26964
rect 17444 26908 17454 26964
rect 28130 26908 28140 26964
rect 28196 26908 29260 26964
rect 29316 26908 29326 26964
rect 12562 26796 12572 26852
rect 12628 26796 13468 26852
rect 13524 26796 13534 26852
rect 17938 26796 17948 26852
rect 18004 26796 19292 26852
rect 19348 26796 26460 26852
rect 26516 26796 29036 26852
rect 29092 26796 30940 26852
rect 30996 26796 32004 26852
rect 31948 26740 32004 26796
rect 22306 26684 22316 26740
rect 22372 26684 22988 26740
rect 23044 26684 23054 26740
rect 31938 26684 31948 26740
rect 32004 26684 34412 26740
rect 34468 26684 34478 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 11218 26460 11228 26516
rect 11284 26460 12908 26516
rect 12964 26460 12974 26516
rect 17714 26460 17724 26516
rect 17780 26460 26236 26516
rect 26292 26460 26302 26516
rect 32498 26460 32508 26516
rect 32564 26460 33404 26516
rect 33460 26460 33470 26516
rect 7522 26348 7532 26404
rect 7588 26348 8316 26404
rect 8372 26348 8382 26404
rect 9538 26348 9548 26404
rect 9604 26348 11116 26404
rect 11172 26348 11182 26404
rect 11330 26348 11340 26404
rect 11396 26348 12684 26404
rect 12740 26348 12750 26404
rect 22530 26348 22540 26404
rect 22596 26348 23212 26404
rect 23268 26348 23278 26404
rect 7970 26236 7980 26292
rect 8036 26236 9660 26292
rect 9716 26236 9726 26292
rect 15250 26236 15260 26292
rect 15316 26236 15932 26292
rect 15988 26236 16492 26292
rect 16548 26236 20860 26292
rect 20916 26236 20926 26292
rect 23426 26236 23436 26292
rect 23492 26236 23884 26292
rect 23940 26236 27356 26292
rect 27412 26236 28364 26292
rect 28420 26236 29932 26292
rect 29988 26236 31164 26292
rect 31220 26236 33964 26292
rect 34020 26236 34030 26292
rect 36530 26236 36540 26292
rect 36596 26236 39004 26292
rect 39060 26236 39070 26292
rect 5618 26124 5628 26180
rect 5684 26124 7868 26180
rect 7924 26124 7934 26180
rect 19954 26124 19964 26180
rect 20020 26124 23772 26180
rect 23828 26124 23996 26180
rect 24052 26124 24062 26180
rect 26674 26124 26684 26180
rect 26740 26124 27692 26180
rect 27748 26124 29148 26180
rect 29204 26124 29214 26180
rect 29474 26124 29484 26180
rect 29540 26124 30380 26180
rect 30436 26124 30446 26180
rect 32834 26124 32844 26180
rect 32900 26124 33292 26180
rect 33348 26124 33358 26180
rect 29586 26012 29596 26068
rect 29652 26012 31612 26068
rect 31668 26012 33516 26068
rect 33572 26012 35308 26068
rect 35364 26012 35374 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 6738 25788 6748 25844
rect 6804 25788 13748 25844
rect 32050 25788 32060 25844
rect 32116 25788 33292 25844
rect 33348 25788 33358 25844
rect 13692 25732 13748 25788
rect 8754 25676 8764 25732
rect 8820 25676 9548 25732
rect 9604 25676 9614 25732
rect 13682 25676 13692 25732
rect 13748 25676 15820 25732
rect 15876 25676 15886 25732
rect 18834 25676 18844 25732
rect 18900 25676 19628 25732
rect 19684 25676 20300 25732
rect 20356 25676 20366 25732
rect 22978 25676 22988 25732
rect 23044 25676 24220 25732
rect 24276 25676 31948 25732
rect 32004 25676 32956 25732
rect 33012 25676 34860 25732
rect 34916 25676 34926 25732
rect 35746 25676 35756 25732
rect 35812 25676 36540 25732
rect 36596 25676 36606 25732
rect 0 25620 800 25648
rect 41200 25620 42000 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 2930 25564 2940 25620
rect 2996 25564 12572 25620
rect 12628 25564 13356 25620
rect 13412 25564 14924 25620
rect 14980 25564 15372 25620
rect 15428 25564 15438 25620
rect 20748 25564 23772 25620
rect 23828 25564 23838 25620
rect 30706 25564 30716 25620
rect 30772 25564 31556 25620
rect 40114 25564 40124 25620
rect 40180 25564 42000 25620
rect 0 25536 800 25564
rect 20748 25508 20804 25564
rect 31500 25508 31556 25564
rect 41200 25536 42000 25564
rect 9762 25452 9772 25508
rect 9828 25452 10444 25508
rect 10500 25452 10510 25508
rect 12002 25452 12012 25508
rect 12068 25452 12460 25508
rect 12516 25452 17052 25508
rect 17108 25452 20804 25508
rect 22866 25452 22876 25508
rect 22932 25452 23660 25508
rect 23716 25452 23726 25508
rect 25218 25452 25228 25508
rect 25284 25452 26796 25508
rect 26852 25452 26862 25508
rect 28802 25452 28812 25508
rect 28868 25452 30828 25508
rect 30884 25452 31276 25508
rect 31332 25452 31342 25508
rect 31490 25452 31500 25508
rect 31556 25452 39004 25508
rect 39060 25452 39070 25508
rect 11218 25340 11228 25396
rect 11284 25340 12124 25396
rect 12180 25340 12190 25396
rect 20626 25340 20636 25396
rect 20692 25340 24444 25396
rect 24500 25340 25452 25396
rect 25508 25340 25518 25396
rect 30258 25340 30268 25396
rect 30324 25340 31164 25396
rect 31220 25340 31230 25396
rect 2818 25228 2828 25284
rect 2884 25228 6636 25284
rect 6692 25228 7644 25284
rect 7700 25228 8652 25284
rect 8708 25228 8718 25284
rect 12786 25228 12796 25284
rect 12852 25228 13468 25284
rect 13524 25228 13534 25284
rect 15698 25228 15708 25284
rect 15764 25228 22540 25284
rect 22596 25228 25564 25284
rect 25620 25228 25630 25284
rect 32498 25228 32508 25284
rect 32564 25228 35756 25284
rect 35812 25228 35822 25284
rect 7970 25116 7980 25172
rect 8036 25116 8540 25172
rect 8596 25116 8606 25172
rect 15810 25116 15820 25172
rect 15876 25116 18732 25172
rect 18788 25116 18798 25172
rect 21970 25116 21980 25172
rect 22036 25116 22428 25172
rect 22484 25116 23324 25172
rect 23380 25116 24444 25172
rect 24500 25116 24510 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 2034 25004 2044 25060
rect 2100 25004 8428 25060
rect 8484 25004 9548 25060
rect 9604 25004 9614 25060
rect 10098 25004 10108 25060
rect 10164 25004 11788 25060
rect 11844 25004 11854 25060
rect 18050 25004 18060 25060
rect 18116 25004 19292 25060
rect 19348 25004 19358 25060
rect 22642 25004 22652 25060
rect 22708 25004 22718 25060
rect 28242 25004 28252 25060
rect 28308 25004 29260 25060
rect 29316 25004 29326 25060
rect 0 24948 800 24976
rect 9548 24948 9604 25004
rect 22652 24948 22708 25004
rect 41200 24948 42000 24976
rect 0 24892 2156 24948
rect 2212 24892 2222 24948
rect 3602 24892 3612 24948
rect 3668 24892 4956 24948
rect 5012 24892 5022 24948
rect 9548 24892 10220 24948
rect 10276 24892 10286 24948
rect 17266 24892 17276 24948
rect 17332 24892 18732 24948
rect 18788 24892 18798 24948
rect 19058 24892 19068 24948
rect 19124 24892 19516 24948
rect 19572 24892 22708 24948
rect 25890 24892 25900 24948
rect 25956 24892 28140 24948
rect 28196 24892 28206 24948
rect 39778 24892 39788 24948
rect 39844 24892 42000 24948
rect 0 24864 800 24892
rect 41200 24864 42000 24892
rect 10658 24780 10668 24836
rect 10724 24780 11340 24836
rect 11396 24780 11406 24836
rect 17388 24780 19740 24836
rect 19796 24780 19806 24836
rect 20514 24780 20524 24836
rect 20580 24780 21532 24836
rect 21588 24780 22988 24836
rect 23044 24780 23054 24836
rect 27234 24780 27244 24836
rect 27300 24780 28476 24836
rect 28532 24780 29372 24836
rect 29428 24780 29438 24836
rect 29586 24780 29596 24836
rect 29652 24780 30492 24836
rect 30548 24780 30558 24836
rect 31714 24780 31724 24836
rect 31780 24780 33068 24836
rect 33124 24780 33134 24836
rect 34626 24780 34636 24836
rect 34692 24780 36204 24836
rect 36260 24780 36270 24836
rect 17388 24724 17444 24780
rect 5394 24668 5404 24724
rect 5460 24668 6524 24724
rect 6580 24668 6860 24724
rect 6916 24668 6926 24724
rect 8978 24668 8988 24724
rect 9044 24668 9996 24724
rect 10052 24668 10062 24724
rect 16370 24668 16380 24724
rect 16436 24668 17388 24724
rect 17444 24668 17454 24724
rect 18610 24668 18620 24724
rect 18676 24668 21644 24724
rect 21700 24668 21710 24724
rect 22082 24668 22092 24724
rect 22148 24668 23996 24724
rect 24052 24668 25228 24724
rect 25284 24668 25900 24724
rect 25956 24668 25966 24724
rect 26674 24668 26684 24724
rect 26740 24668 28588 24724
rect 28644 24668 28654 24724
rect 33170 24668 33180 24724
rect 33236 24668 34188 24724
rect 34244 24668 36316 24724
rect 36372 24668 36382 24724
rect 16818 24556 16828 24612
rect 16884 24556 17500 24612
rect 17556 24556 17566 24612
rect 19730 24556 19740 24612
rect 19796 24556 20300 24612
rect 20356 24556 20366 24612
rect 23762 24556 23772 24612
rect 23828 24556 25004 24612
rect 25060 24556 25070 24612
rect 34402 24556 34412 24612
rect 34468 24556 35644 24612
rect 35700 24556 35710 24612
rect 9986 24444 9996 24500
rect 10052 24444 11228 24500
rect 11284 24444 11294 24500
rect 32050 24444 32060 24500
rect 32116 24444 33516 24500
rect 33572 24444 35420 24500
rect 35476 24444 35486 24500
rect 0 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 0 24220 1708 24276
rect 1764 24220 2492 24276
rect 2548 24220 2558 24276
rect 0 24192 800 24220
rect 7074 23996 7084 24052
rect 7140 23996 8540 24052
rect 8596 23996 8606 24052
rect 13234 23996 13244 24052
rect 13300 23996 14476 24052
rect 14532 23996 14542 24052
rect 2258 23884 2268 23940
rect 2324 23884 2334 23940
rect 7186 23884 7196 23940
rect 7252 23884 10556 23940
rect 10612 23884 11564 23940
rect 11620 23884 11630 23940
rect 20626 23884 20636 23940
rect 20692 23884 20972 23940
rect 21028 23884 21038 23940
rect 21634 23884 21644 23940
rect 21700 23884 22428 23940
rect 22484 23884 22494 23940
rect 23202 23884 23212 23940
rect 23268 23884 23996 23940
rect 24052 23884 24062 23940
rect 28354 23884 28364 23940
rect 28420 23884 30380 23940
rect 30436 23884 30446 23940
rect 32386 23884 32396 23940
rect 32452 23884 33068 23940
rect 33124 23884 34300 23940
rect 34356 23884 35420 23940
rect 35476 23884 35868 23940
rect 35924 23884 35934 23940
rect 38612 23884 39004 23940
rect 39060 23884 39070 23940
rect 2268 23828 2324 23884
rect 2268 23772 9436 23828
rect 9492 23772 10444 23828
rect 10500 23772 12012 23828
rect 12068 23772 13468 23828
rect 13524 23772 13534 23828
rect 18050 23772 18060 23828
rect 18116 23772 18732 23828
rect 18788 23772 19516 23828
rect 19572 23772 19582 23828
rect 20738 23772 20748 23828
rect 20804 23772 22092 23828
rect 22148 23772 22652 23828
rect 22708 23772 24332 23828
rect 24388 23772 24398 23828
rect 26002 23772 26012 23828
rect 26068 23772 26684 23828
rect 26740 23772 26750 23828
rect 28242 23772 28252 23828
rect 28308 23772 30492 23828
rect 30548 23772 30558 23828
rect 38612 23716 38668 23884
rect 8082 23660 8092 23716
rect 8148 23660 8764 23716
rect 8820 23660 9772 23716
rect 9828 23660 9838 23716
rect 13682 23660 13692 23716
rect 13748 23660 15148 23716
rect 15204 23660 15214 23716
rect 18610 23660 18620 23716
rect 18676 23660 19404 23716
rect 19460 23660 19470 23716
rect 28130 23660 28140 23716
rect 28196 23660 30268 23716
rect 30324 23660 38668 23716
rect 0 23604 800 23632
rect 41200 23604 42000 23632
rect 0 23548 1708 23604
rect 1764 23548 2716 23604
rect 2772 23548 2782 23604
rect 16370 23548 16380 23604
rect 16436 23548 17276 23604
rect 17332 23548 17342 23604
rect 29474 23548 29484 23604
rect 29540 23548 30604 23604
rect 30660 23548 36764 23604
rect 36820 23548 38332 23604
rect 38388 23548 38398 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 9538 23436 9548 23492
rect 9604 23436 10220 23492
rect 10276 23436 10286 23492
rect 11666 23436 11676 23492
rect 11732 23436 19628 23492
rect 19684 23436 19694 23492
rect 20524 23436 21980 23492
rect 22036 23436 22046 23492
rect 20524 23380 20580 23436
rect 2818 23324 2828 23380
rect 2884 23324 3388 23380
rect 3444 23324 16828 23380
rect 16884 23324 16894 23380
rect 18386 23324 18396 23380
rect 18452 23324 19292 23380
rect 19348 23324 19358 23380
rect 19954 23324 19964 23380
rect 20020 23324 20580 23380
rect 20738 23324 20748 23380
rect 20804 23324 21084 23380
rect 21140 23324 21150 23380
rect 21858 23324 21868 23380
rect 21924 23324 22876 23380
rect 22932 23324 22942 23380
rect 29698 23324 29708 23380
rect 29764 23324 32172 23380
rect 32228 23324 33292 23380
rect 33348 23324 33358 23380
rect 8082 23212 8092 23268
rect 8148 23212 8316 23268
rect 8372 23212 9660 23268
rect 9716 23212 9726 23268
rect 10322 23212 10332 23268
rect 10388 23212 11116 23268
rect 11172 23212 12124 23268
rect 12180 23212 12190 23268
rect 17490 23212 17500 23268
rect 17556 23212 17566 23268
rect 19618 23212 19628 23268
rect 19684 23212 20412 23268
rect 20468 23212 27692 23268
rect 27748 23212 27758 23268
rect 34066 23212 34076 23268
rect 34132 23212 34636 23268
rect 34692 23212 34702 23268
rect 17500 23156 17556 23212
rect 7298 23100 7308 23156
rect 7364 23100 9548 23156
rect 9604 23100 9614 23156
rect 15362 23100 15372 23156
rect 15428 23100 17556 23156
rect 17714 23100 17724 23156
rect 17780 23100 18396 23156
rect 18452 23100 18462 23156
rect 20962 23100 20972 23156
rect 21028 23100 21644 23156
rect 21700 23100 21710 23156
rect 24546 23100 24556 23156
rect 24612 23100 26460 23156
rect 26516 23100 26526 23156
rect 1922 22988 1932 23044
rect 1988 22988 1998 23044
rect 19282 22988 19292 23044
rect 19348 22988 19964 23044
rect 20020 22988 20030 23044
rect 21186 22988 21196 23044
rect 21252 22988 21868 23044
rect 21924 22988 21934 23044
rect 24210 22988 24220 23044
rect 24276 22988 24780 23044
rect 24836 22988 25676 23044
rect 25732 22988 25742 23044
rect 26226 22988 26236 23044
rect 26292 22988 26796 23044
rect 26852 22988 27692 23044
rect 27748 22988 28700 23044
rect 28756 22988 28766 23044
rect 29922 22988 29932 23044
rect 29988 22988 31164 23044
rect 31220 22988 31230 23044
rect 38546 22988 38556 23044
rect 0 22932 800 22960
rect 1932 22932 1988 22988
rect 21868 22932 21924 22988
rect 38612 22932 38668 23044
rect 41200 22932 42000 22960
rect 0 22876 1988 22932
rect 9762 22876 9772 22932
rect 9828 22876 11340 22932
rect 11396 22876 11406 22932
rect 16258 22876 16268 22932
rect 16324 22876 18060 22932
rect 18116 22876 18126 22932
rect 21868 22876 25900 22932
rect 25956 22876 25966 22932
rect 27234 22876 27244 22932
rect 27300 22876 29036 22932
rect 29092 22876 29102 22932
rect 38612 22876 40236 22932
rect 40292 22876 42000 22932
rect 0 22848 800 22876
rect 41200 22848 42000 22876
rect 8642 22764 8652 22820
rect 8708 22764 9212 22820
rect 9268 22764 9278 22820
rect 21746 22764 21756 22820
rect 21812 22764 22876 22820
rect 22932 22764 22942 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 8418 22540 8428 22596
rect 8484 22540 9324 22596
rect 9380 22540 9390 22596
rect 21858 22540 21868 22596
rect 21924 22540 22204 22596
rect 22260 22540 22270 22596
rect 28578 22540 28588 22596
rect 28644 22540 29484 22596
rect 29540 22540 29550 22596
rect 5058 22428 5068 22484
rect 5124 22428 5740 22484
rect 5796 22428 5806 22484
rect 7522 22428 7532 22484
rect 7588 22428 7980 22484
rect 8036 22428 8652 22484
rect 8708 22428 8718 22484
rect 12898 22428 12908 22484
rect 12964 22428 13692 22484
rect 13748 22428 15932 22484
rect 15988 22428 23100 22484
rect 23156 22428 23166 22484
rect 28466 22428 28476 22484
rect 28532 22428 30156 22484
rect 30212 22428 31388 22484
rect 31444 22428 31454 22484
rect 31602 22428 31612 22484
rect 31668 22428 32844 22484
rect 32900 22428 32910 22484
rect 35074 22428 35084 22484
rect 35140 22428 35868 22484
rect 35924 22428 35934 22484
rect 6402 22316 6412 22372
rect 6468 22316 8764 22372
rect 8820 22316 10220 22372
rect 10276 22316 10286 22372
rect 11218 22316 11228 22372
rect 11284 22316 12684 22372
rect 12740 22316 12750 22372
rect 24434 22316 24444 22372
rect 24500 22316 25788 22372
rect 25844 22316 25854 22372
rect 32946 22316 32956 22372
rect 33012 22316 33516 22372
rect 33572 22316 34972 22372
rect 35028 22316 35038 22372
rect 0 22260 800 22288
rect 41200 22260 42000 22288
rect 0 22204 1932 22260
rect 1988 22204 3276 22260
rect 3332 22204 3342 22260
rect 8418 22204 8428 22260
rect 8484 22204 11900 22260
rect 11956 22204 11966 22260
rect 16594 22204 16604 22260
rect 16660 22204 17164 22260
rect 17220 22204 17230 22260
rect 32274 22204 32284 22260
rect 32340 22204 33404 22260
rect 33460 22204 33852 22260
rect 33908 22204 35420 22260
rect 35476 22204 35486 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 0 22176 800 22204
rect 41200 22176 42000 22204
rect 1586 22092 1596 22148
rect 1652 22092 2828 22148
rect 2884 22092 5628 22148
rect 5684 22092 6188 22148
rect 6244 22092 6524 22148
rect 6580 22092 6590 22148
rect 8866 22092 8876 22148
rect 8932 22092 10444 22148
rect 10500 22092 10510 22148
rect 10882 22092 10892 22148
rect 10948 22092 13468 22148
rect 13524 22092 13534 22148
rect 14690 22092 14700 22148
rect 14756 22092 17388 22148
rect 17444 22092 17454 22148
rect 18162 22092 18172 22148
rect 18228 22092 18956 22148
rect 19012 22092 19022 22148
rect 19954 22092 19964 22148
rect 20020 22092 20524 22148
rect 20580 22092 20748 22148
rect 20804 22092 22204 22148
rect 22260 22092 22270 22148
rect 25442 22092 25452 22148
rect 25508 22092 27468 22148
rect 27524 22092 39900 22148
rect 39956 22092 39966 22148
rect 8082 21980 8092 22036
rect 8148 21980 9436 22036
rect 9492 21980 9502 22036
rect 17938 21980 17948 22036
rect 18004 21980 18732 22036
rect 18788 21980 19292 22036
rect 19348 21980 19358 22036
rect 20290 21980 20300 22036
rect 20356 21980 21532 22036
rect 21588 21980 21598 22036
rect 33068 21980 33180 22036
rect 33236 21980 33246 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 9762 21868 9772 21924
rect 9828 21868 10220 21924
rect 10276 21868 10286 21924
rect 10434 21868 10444 21924
rect 10500 21868 11340 21924
rect 11396 21868 11406 21924
rect 20300 21812 20356 21980
rect 2370 21756 2380 21812
rect 2436 21756 4732 21812
rect 4788 21756 4798 21812
rect 5730 21756 5740 21812
rect 5796 21756 6748 21812
rect 6804 21756 6814 21812
rect 12898 21756 12908 21812
rect 12964 21756 14028 21812
rect 14084 21756 14094 21812
rect 17490 21756 17500 21812
rect 17556 21756 17724 21812
rect 17780 21756 19292 21812
rect 19348 21756 20356 21812
rect 21410 21756 21420 21812
rect 21476 21756 25340 21812
rect 25396 21756 25406 21812
rect 30034 21756 30044 21812
rect 30100 21756 30940 21812
rect 30996 21756 31006 21812
rect 31490 21756 31500 21812
rect 31556 21756 32732 21812
rect 32788 21756 32798 21812
rect 33068 21700 33124 21980
rect 33282 21868 33292 21924
rect 33348 21868 33358 21924
rect 33292 21812 33348 21868
rect 33292 21756 33740 21812
rect 33796 21756 33806 21812
rect 3826 21644 3836 21700
rect 3892 21644 6188 21700
rect 6244 21644 6636 21700
rect 6692 21644 6702 21700
rect 11442 21644 11452 21700
rect 11508 21644 12572 21700
rect 12628 21644 12638 21700
rect 16482 21644 16492 21700
rect 16548 21644 16828 21700
rect 16884 21644 17948 21700
rect 18004 21644 18014 21700
rect 20738 21644 20748 21700
rect 20804 21644 22428 21700
rect 22484 21644 23660 21700
rect 23716 21644 23726 21700
rect 26562 21644 26572 21700
rect 26628 21644 27580 21700
rect 27636 21644 27646 21700
rect 28466 21644 28476 21700
rect 28532 21644 29260 21700
rect 29316 21644 29326 21700
rect 33068 21644 33628 21700
rect 33684 21644 33694 21700
rect 33842 21644 33852 21700
rect 33908 21644 34636 21700
rect 34692 21644 34702 21700
rect 0 21588 800 21616
rect 41200 21588 42000 21616
rect 0 21532 2156 21588
rect 2212 21532 2222 21588
rect 4050 21532 4060 21588
rect 4116 21532 18508 21588
rect 18564 21532 18574 21588
rect 0 21504 800 21532
rect 17042 21420 17052 21476
rect 17108 21420 18284 21476
rect 18340 21420 18350 21476
rect 26852 21364 26908 21588
rect 26964 21532 26974 21588
rect 28354 21532 28364 21588
rect 28420 21532 29708 21588
rect 29764 21532 29774 21588
rect 30258 21532 30268 21588
rect 30324 21532 30828 21588
rect 30884 21532 30894 21588
rect 32498 21532 32508 21588
rect 32564 21532 33964 21588
rect 34020 21532 34030 21588
rect 37986 21532 37996 21588
rect 38052 21532 39116 21588
rect 39172 21532 39182 21588
rect 39554 21532 39564 21588
rect 39620 21532 42000 21588
rect 32508 21476 32564 21532
rect 41200 21504 42000 21532
rect 31836 21420 32564 21476
rect 31836 21364 31892 21420
rect 13458 21308 13468 21364
rect 13524 21308 14924 21364
rect 14980 21308 14990 21364
rect 24210 21308 24220 21364
rect 24276 21308 26908 21364
rect 31826 21308 31836 21364
rect 31892 21308 31902 21364
rect 33282 21308 33292 21364
rect 33348 21308 35084 21364
rect 35140 21308 35150 21364
rect 33292 21252 33348 21308
rect 17602 21196 17612 21252
rect 17668 21196 18284 21252
rect 18340 21196 19852 21252
rect 19908 21196 19918 21252
rect 23538 21196 23548 21252
rect 23604 21196 25452 21252
rect 25508 21196 25518 21252
rect 28914 21196 28924 21252
rect 28980 21196 33348 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 18610 21084 18620 21140
rect 18676 21084 18686 21140
rect 24658 21084 24668 21140
rect 24724 21084 26012 21140
rect 26068 21084 26078 21140
rect 18620 21028 18676 21084
rect 4498 20972 4508 21028
rect 4564 20972 8204 21028
rect 8260 20972 8270 21028
rect 14466 20972 14476 21028
rect 14532 20972 15932 21028
rect 15988 20972 18060 21028
rect 18116 20972 18676 21028
rect 22194 20972 22204 21028
rect 22260 20972 23324 21028
rect 23380 20972 26684 21028
rect 26740 20972 26750 21028
rect 29250 20972 29260 21028
rect 29316 20972 30604 21028
rect 30660 20972 30670 21028
rect 33628 20972 35420 21028
rect 35476 20972 37996 21028
rect 38052 20972 38062 21028
rect 0 20916 800 20944
rect 33628 20916 33684 20972
rect 41200 20916 42000 20944
rect 0 20860 1708 20916
rect 1764 20860 3724 20916
rect 3780 20860 3790 20916
rect 15698 20860 15708 20916
rect 15764 20860 18396 20916
rect 18452 20860 18462 20916
rect 20178 20860 20188 20916
rect 20244 20860 20524 20916
rect 20580 20860 20590 20916
rect 22866 20860 22876 20916
rect 22932 20860 24220 20916
rect 24276 20860 24286 20916
rect 31714 20860 31724 20916
rect 31780 20860 33628 20916
rect 33684 20860 33694 20916
rect 34402 20860 34412 20916
rect 34468 20860 35532 20916
rect 35588 20860 35598 20916
rect 40114 20860 40124 20916
rect 40180 20860 42000 20916
rect 0 20832 800 20860
rect 41200 20832 42000 20860
rect 4274 20748 4284 20804
rect 4340 20748 5964 20804
rect 6020 20748 6030 20804
rect 6178 20748 6188 20804
rect 6244 20748 6524 20804
rect 6580 20748 7196 20804
rect 7252 20748 7262 20804
rect 9650 20748 9660 20804
rect 9716 20748 10108 20804
rect 10164 20748 10174 20804
rect 12338 20748 12348 20804
rect 12404 20748 13468 20804
rect 13524 20748 13534 20804
rect 17042 20748 17052 20804
rect 17108 20748 17724 20804
rect 17780 20748 18620 20804
rect 18676 20748 18686 20804
rect 22642 20748 22652 20804
rect 22708 20748 23996 20804
rect 24052 20748 24062 20804
rect 27682 20748 27692 20804
rect 27748 20748 30156 20804
rect 30212 20748 30222 20804
rect 32834 20748 32844 20804
rect 32900 20748 35084 20804
rect 35140 20748 35150 20804
rect 4732 20692 4788 20748
rect 4722 20636 4732 20692
rect 4788 20636 4798 20692
rect 6626 20636 6636 20692
rect 6692 20636 7420 20692
rect 7476 20636 8428 20692
rect 8484 20636 9212 20692
rect 9268 20636 9278 20692
rect 14242 20636 14252 20692
rect 14308 20636 18844 20692
rect 18900 20636 18910 20692
rect 19842 20636 19852 20692
rect 19908 20636 20860 20692
rect 20916 20636 20926 20692
rect 21746 20636 21756 20692
rect 21812 20636 23772 20692
rect 23828 20636 23838 20692
rect 33730 20636 33740 20692
rect 33796 20636 35196 20692
rect 35252 20636 35262 20692
rect 18844 20580 18900 20636
rect 16034 20524 16044 20580
rect 16100 20524 17836 20580
rect 17892 20524 17902 20580
rect 18844 20524 22092 20580
rect 22148 20524 22158 20580
rect 23650 20524 23660 20580
rect 23716 20524 24444 20580
rect 24500 20524 24510 20580
rect 25564 20524 28588 20580
rect 28644 20524 29260 20580
rect 29316 20524 29326 20580
rect 31266 20524 31276 20580
rect 31332 20524 32060 20580
rect 32116 20524 32620 20580
rect 32676 20524 32686 20580
rect 34514 20524 34524 20580
rect 34580 20524 34972 20580
rect 35028 20524 36092 20580
rect 36148 20524 36158 20580
rect 16370 20412 16380 20468
rect 16436 20412 17724 20468
rect 17780 20412 17790 20468
rect 17938 20412 17948 20468
rect 18004 20412 18396 20468
rect 18452 20412 18462 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 25564 20356 25620 20524
rect 25778 20412 25788 20468
rect 25844 20412 39004 20468
rect 39060 20412 39070 20468
rect 6066 20300 6076 20356
rect 6132 20300 6412 20356
rect 6468 20300 6478 20356
rect 7634 20300 7644 20356
rect 7700 20300 8876 20356
rect 8932 20300 10220 20356
rect 10276 20300 10286 20356
rect 17826 20300 17836 20356
rect 17892 20300 18004 20356
rect 22978 20300 22988 20356
rect 23044 20300 24220 20356
rect 24276 20300 25620 20356
rect 0 20244 800 20272
rect 0 20188 2604 20244
rect 2660 20188 3612 20244
rect 3668 20188 3678 20244
rect 10322 20188 10332 20244
rect 10388 20188 10780 20244
rect 10836 20188 10846 20244
rect 11732 20188 14028 20244
rect 14084 20188 14094 20244
rect 17042 20188 17052 20244
rect 17108 20188 17724 20244
rect 17780 20188 17790 20244
rect 0 20160 800 20188
rect 2258 20076 2268 20132
rect 2324 20076 3388 20132
rect 4162 20076 4172 20132
rect 4228 20076 5180 20132
rect 5236 20076 5628 20132
rect 5684 20076 6972 20132
rect 7028 20076 7038 20132
rect 8306 20076 8316 20132
rect 8372 20076 9548 20132
rect 9604 20076 9614 20132
rect 10882 20076 10892 20132
rect 10948 20076 10958 20132
rect 3332 20020 3388 20076
rect 10892 20020 10948 20076
rect 11732 20020 11788 20188
rect 17948 20132 18004 20300
rect 41200 20244 42000 20272
rect 23986 20188 23996 20244
rect 24052 20188 25228 20244
rect 25284 20188 25294 20244
rect 39666 20188 39676 20244
rect 39732 20188 40236 20244
rect 40292 20188 42000 20244
rect 41200 20160 42000 20188
rect 15810 20076 15820 20132
rect 15876 20076 18004 20132
rect 25442 20076 25452 20132
rect 25508 20076 26236 20132
rect 26292 20076 26302 20132
rect 26562 20076 26572 20132
rect 26628 20076 29148 20132
rect 29204 20076 29214 20132
rect 34178 20076 34188 20132
rect 34244 20076 38444 20132
rect 38500 20076 38510 20132
rect 38612 20076 39228 20132
rect 39284 20076 39294 20132
rect 3332 19964 7644 20020
rect 7700 19964 7710 20020
rect 7858 19964 7868 20020
rect 7924 19964 8428 20020
rect 8484 19964 8494 20020
rect 10434 19964 10444 20020
rect 10500 19964 11788 20020
rect 14578 19964 14588 20020
rect 14644 19964 16716 20020
rect 16772 19964 18732 20020
rect 18788 19964 18798 20020
rect 24770 19964 24780 20020
rect 24836 19964 26684 20020
rect 26740 19964 26750 20020
rect 29250 19964 29260 20020
rect 29316 19964 30380 20020
rect 30436 19964 30446 20020
rect 31490 19964 31500 20020
rect 31556 19964 31948 20020
rect 32004 19964 32284 20020
rect 32340 19964 32350 20020
rect 38612 19908 38668 20076
rect 7970 19852 7980 19908
rect 8036 19852 10892 19908
rect 10948 19852 10958 19908
rect 17826 19852 17836 19908
rect 17892 19852 22764 19908
rect 22820 19852 22830 19908
rect 26226 19852 26236 19908
rect 26292 19852 27244 19908
rect 27300 19852 38668 19908
rect 3154 19740 3164 19796
rect 3220 19740 14252 19796
rect 14308 19740 15036 19796
rect 7634 19628 7644 19684
rect 7700 19628 12236 19684
rect 12292 19628 12302 19684
rect 0 19572 800 19600
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 0 19516 1932 19572
rect 1988 19516 1998 19572
rect 0 19488 800 19516
rect 7522 19404 7532 19460
rect 7588 19404 8540 19460
rect 8596 19404 8606 19460
rect 15092 19404 15148 19796
rect 24546 19740 24556 19796
rect 24612 19740 26572 19796
rect 26628 19740 26638 19796
rect 29922 19740 29932 19796
rect 29988 19740 31276 19796
rect 31332 19740 32508 19796
rect 32564 19740 32574 19796
rect 24098 19628 24108 19684
rect 24164 19628 26460 19684
rect 26516 19628 26526 19684
rect 29698 19628 29708 19684
rect 29764 19628 31052 19684
rect 31108 19628 31118 19684
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 24658 19516 24668 19572
rect 24724 19516 33628 19572
rect 33684 19516 33694 19572
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 33628 19460 33684 19516
rect 41200 19488 42000 19516
rect 15204 19404 15820 19460
rect 15876 19404 15886 19460
rect 24322 19404 24332 19460
rect 24388 19404 25340 19460
rect 25396 19404 26124 19460
rect 26180 19404 26190 19460
rect 33628 19404 35532 19460
rect 35588 19404 35598 19460
rect 4498 19292 4508 19348
rect 4564 19292 8764 19348
rect 8820 19292 8830 19348
rect 12450 19292 12460 19348
rect 12516 19292 13916 19348
rect 13972 19292 15036 19348
rect 15092 19292 15102 19348
rect 15362 19292 15372 19348
rect 15428 19292 16044 19348
rect 16100 19292 16110 19348
rect 20402 19292 20412 19348
rect 20468 19292 22204 19348
rect 22260 19292 22270 19348
rect 39890 19292 39900 19348
rect 39956 19292 39966 19348
rect 39900 19236 39956 19292
rect 2930 19180 2940 19236
rect 2996 19180 5740 19236
rect 5796 19180 6300 19236
rect 6356 19180 6366 19236
rect 10882 19180 10892 19236
rect 10948 19180 11284 19236
rect 12898 19180 12908 19236
rect 12964 19180 13468 19236
rect 13524 19180 13534 19236
rect 16818 19180 16828 19236
rect 16884 19180 17724 19236
rect 17780 19180 17790 19236
rect 24098 19180 24108 19236
rect 24164 19180 25676 19236
rect 25732 19180 25900 19236
rect 25956 19180 25966 19236
rect 28466 19180 28476 19236
rect 28532 19180 28542 19236
rect 30146 19180 30156 19236
rect 30212 19180 30716 19236
rect 30772 19180 39956 19236
rect 2034 19068 2044 19124
rect 2100 19068 2110 19124
rect 3602 19068 3612 19124
rect 3668 19068 10668 19124
rect 10724 19068 11004 19124
rect 11060 19068 11070 19124
rect 0 18900 800 18928
rect 2044 18900 2100 19068
rect 11228 19012 11284 19180
rect 12674 19068 12684 19124
rect 12740 19068 13916 19124
rect 13972 19068 14588 19124
rect 14644 19068 14654 19124
rect 19506 19068 19516 19124
rect 19572 19068 21420 19124
rect 21476 19068 21486 19124
rect 24882 19068 24892 19124
rect 24948 19068 26236 19124
rect 26292 19068 26302 19124
rect 28476 19012 28532 19180
rect 31042 19068 31052 19124
rect 31108 19068 32620 19124
rect 32676 19068 34076 19124
rect 34132 19068 34142 19124
rect 3154 18956 3164 19012
rect 3220 18956 4172 19012
rect 4228 18956 4238 19012
rect 8754 18956 8764 19012
rect 8820 18956 9324 19012
rect 9380 18956 10220 19012
rect 10276 18956 17724 19012
rect 17780 18956 17790 19012
rect 20290 18956 20300 19012
rect 20356 18956 21308 19012
rect 21364 18956 21374 19012
rect 28476 18956 39900 19012
rect 39956 18956 39966 19012
rect 41200 18900 42000 18928
rect 0 18844 2100 18900
rect 12898 18844 12908 18900
rect 12964 18844 13692 18900
rect 13748 18844 14700 18900
rect 14756 18844 14766 18900
rect 31154 18844 31164 18900
rect 31220 18844 31500 18900
rect 31556 18844 31566 18900
rect 32722 18844 32732 18900
rect 32788 18844 33516 18900
rect 33572 18844 33582 18900
rect 39666 18844 39676 18900
rect 39732 18844 40236 18900
rect 40292 18844 42000 18900
rect 0 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 41200 18816 42000 18844
rect 10210 18732 10220 18788
rect 10276 18732 10780 18788
rect 10836 18732 11676 18788
rect 11732 18732 11742 18788
rect 13346 18732 13356 18788
rect 13412 18732 14028 18788
rect 14084 18732 14094 18788
rect 6178 18620 6188 18676
rect 6244 18620 6860 18676
rect 6916 18620 6926 18676
rect 2706 18508 2716 18564
rect 2772 18508 3724 18564
rect 3780 18508 3790 18564
rect 6962 18508 6972 18564
rect 7028 18508 7532 18564
rect 7588 18508 9772 18564
rect 9828 18508 19180 18564
rect 19236 18508 19246 18564
rect 19180 18452 19236 18508
rect 2146 18396 2156 18452
rect 2212 18396 6524 18452
rect 6580 18396 6590 18452
rect 10770 18396 10780 18452
rect 10836 18396 11452 18452
rect 11508 18396 11518 18452
rect 12002 18396 12012 18452
rect 12068 18396 12796 18452
rect 12852 18396 12862 18452
rect 15250 18396 15260 18452
rect 15316 18396 16268 18452
rect 16324 18396 16334 18452
rect 16482 18396 16492 18452
rect 16548 18396 17836 18452
rect 17892 18396 17902 18452
rect 19180 18396 21644 18452
rect 21700 18396 21710 18452
rect 25778 18396 25788 18452
rect 25844 18396 26796 18452
rect 26852 18396 26862 18452
rect 11452 18340 11508 18396
rect 2594 18284 2604 18340
rect 2660 18284 4620 18340
rect 4676 18284 4686 18340
rect 11452 18284 12572 18340
rect 12628 18284 12638 18340
rect 16370 18284 16380 18340
rect 16436 18284 16828 18340
rect 16884 18284 18060 18340
rect 18116 18284 18126 18340
rect 21410 18284 21420 18340
rect 21476 18284 21980 18340
rect 22036 18284 22988 18340
rect 23044 18284 23054 18340
rect 26338 18284 26348 18340
rect 26404 18284 27356 18340
rect 27412 18284 27422 18340
rect 27570 18284 27580 18340
rect 27636 18284 29148 18340
rect 29204 18284 29214 18340
rect 31714 18284 31724 18340
rect 31780 18284 32172 18340
rect 32228 18284 33740 18340
rect 33796 18284 34748 18340
rect 34804 18284 35532 18340
rect 35588 18284 35598 18340
rect 0 18228 800 18256
rect 0 18172 2100 18228
rect 2258 18172 2268 18228
rect 2324 18172 10836 18228
rect 11330 18172 11340 18228
rect 11396 18172 14364 18228
rect 14420 18172 14430 18228
rect 19394 18172 19404 18228
rect 19460 18172 20412 18228
rect 20468 18172 23772 18228
rect 23828 18172 23838 18228
rect 33842 18172 33852 18228
rect 33908 18172 34524 18228
rect 34580 18172 34590 18228
rect 0 18144 800 18172
rect 2044 18116 2100 18172
rect 10780 18116 10836 18172
rect 2044 18060 3388 18116
rect 3444 18060 3454 18116
rect 10780 18060 12236 18116
rect 12292 18060 12796 18116
rect 12852 18060 12862 18116
rect 18946 18060 18956 18116
rect 19012 18060 19964 18116
rect 20020 18060 21644 18116
rect 21700 18060 24556 18116
rect 24612 18060 24622 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 11442 17948 11452 18004
rect 11508 17948 13468 18004
rect 13524 17948 13534 18004
rect 21186 17948 21196 18004
rect 21252 17948 22428 18004
rect 22484 17948 23212 18004
rect 23268 17948 23660 18004
rect 23716 17948 24108 18004
rect 24164 17948 24174 18004
rect 13010 17836 13020 17892
rect 13076 17836 14252 17892
rect 14308 17836 14318 17892
rect 14476 17836 16380 17892
rect 16436 17836 16446 17892
rect 19730 17836 19740 17892
rect 19796 17836 20412 17892
rect 20468 17836 21308 17892
rect 21364 17836 21374 17892
rect 21532 17836 26348 17892
rect 26404 17836 26414 17892
rect 10994 17724 11004 17780
rect 11060 17724 11452 17780
rect 11508 17724 11518 17780
rect 13458 17724 13468 17780
rect 13524 17724 14140 17780
rect 14196 17724 14206 17780
rect 14476 17668 14532 17836
rect 21532 17780 21588 17836
rect 14690 17724 14700 17780
rect 14756 17724 16604 17780
rect 16660 17724 17164 17780
rect 17220 17724 17230 17780
rect 18386 17724 18396 17780
rect 18452 17724 19292 17780
rect 19348 17724 19852 17780
rect 19908 17724 19918 17780
rect 20738 17724 20748 17780
rect 20804 17724 21588 17780
rect 25890 17724 25900 17780
rect 25956 17724 29372 17780
rect 29428 17724 30044 17780
rect 30100 17724 34636 17780
rect 34692 17724 35980 17780
rect 36036 17724 36046 17780
rect 8530 17612 8540 17668
rect 8596 17612 10332 17668
rect 10388 17612 10398 17668
rect 10658 17612 10668 17668
rect 10724 17612 11788 17668
rect 11844 17612 11854 17668
rect 12012 17612 14532 17668
rect 14588 17612 15372 17668
rect 15428 17612 15438 17668
rect 18162 17612 18172 17668
rect 18228 17612 21868 17668
rect 21924 17612 21934 17668
rect 22754 17612 22764 17668
rect 22820 17612 25452 17668
rect 25508 17612 25518 17668
rect 29250 17612 29260 17668
rect 29316 17612 29708 17668
rect 29764 17612 31388 17668
rect 31444 17612 31454 17668
rect 0 17556 800 17584
rect 12012 17556 12068 17612
rect 14588 17556 14644 17612
rect 0 17500 1708 17556
rect 1764 17500 1774 17556
rect 3714 17500 3724 17556
rect 3780 17500 12068 17556
rect 12674 17500 12684 17556
rect 12740 17500 13468 17556
rect 13524 17500 13534 17556
rect 14354 17500 14364 17556
rect 14420 17500 14644 17556
rect 14914 17500 14924 17556
rect 14980 17500 21532 17556
rect 21588 17500 21598 17556
rect 34962 17500 34972 17556
rect 35028 17500 35532 17556
rect 35588 17500 35598 17556
rect 0 17472 800 17500
rect 14924 17444 14980 17500
rect 2594 17388 2604 17444
rect 2660 17388 4060 17444
rect 4116 17388 4126 17444
rect 5058 17388 5068 17444
rect 5124 17388 9548 17444
rect 9604 17388 9614 17444
rect 14018 17388 14028 17444
rect 14084 17388 14980 17444
rect 15362 17388 15372 17444
rect 15428 17388 20748 17444
rect 20804 17388 20814 17444
rect 25218 17388 25228 17444
rect 25284 17388 26516 17444
rect 26674 17388 26684 17444
rect 26740 17388 28028 17444
rect 28084 17388 28094 17444
rect 32834 17388 32844 17444
rect 32900 17388 34524 17444
rect 34580 17388 34590 17444
rect 26460 17332 26516 17388
rect 8530 17276 8540 17332
rect 8596 17276 9100 17332
rect 9156 17276 12012 17332
rect 12068 17276 17052 17332
rect 17108 17276 17118 17332
rect 21522 17276 21532 17332
rect 21588 17276 23100 17332
rect 23156 17276 25732 17332
rect 26460 17276 28476 17332
rect 28532 17276 29820 17332
rect 29876 17276 29886 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 25676 17108 25732 17276
rect 2930 17052 2940 17108
rect 2996 17052 9996 17108
rect 10052 17052 10444 17108
rect 10500 17052 10780 17108
rect 10836 17052 10846 17108
rect 11890 17052 11900 17108
rect 11956 17052 13244 17108
rect 13300 17052 13310 17108
rect 22978 17052 22988 17108
rect 23044 17052 25228 17108
rect 25284 17052 25294 17108
rect 25676 17052 32060 17108
rect 32116 17052 32126 17108
rect 10098 16940 10108 16996
rect 10164 16940 14252 16996
rect 14308 16940 14812 16996
rect 14868 16940 17388 16996
rect 17444 16940 17454 16996
rect 24546 16940 24556 16996
rect 24612 16940 26124 16996
rect 26180 16940 26572 16996
rect 26628 16940 26638 16996
rect 26786 16940 26796 16996
rect 26852 16940 27804 16996
rect 27860 16940 28476 16996
rect 28532 16940 28542 16996
rect 29810 16940 29820 16996
rect 29876 16940 33292 16996
rect 33348 16940 33358 16996
rect 34178 16940 34188 16996
rect 34244 16940 37212 16996
rect 37268 16940 37278 16996
rect 0 16884 800 16912
rect 41200 16884 42000 16912
rect 0 16828 2604 16884
rect 2660 16828 2670 16884
rect 12450 16828 12460 16884
rect 12516 16828 13916 16884
rect 13972 16828 13982 16884
rect 15922 16828 15932 16884
rect 15988 16828 17276 16884
rect 17332 16828 17342 16884
rect 19954 16828 19964 16884
rect 20020 16828 21980 16884
rect 22036 16828 22046 16884
rect 22418 16828 22428 16884
rect 22484 16828 28700 16884
rect 28756 16828 28766 16884
rect 31378 16828 31388 16884
rect 31444 16828 33628 16884
rect 33684 16828 34860 16884
rect 34916 16828 34926 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 0 16800 800 16828
rect 41200 16800 42000 16828
rect 7298 16716 7308 16772
rect 7364 16716 8988 16772
rect 9044 16716 9054 16772
rect 15250 16716 15260 16772
rect 15316 16716 15596 16772
rect 15652 16716 16268 16772
rect 16324 16716 16828 16772
rect 16884 16716 17612 16772
rect 17668 16716 17678 16772
rect 18386 16716 18396 16772
rect 18452 16716 19628 16772
rect 19684 16716 19694 16772
rect 25890 16716 25900 16772
rect 25956 16716 27020 16772
rect 27076 16716 27086 16772
rect 10882 16604 10892 16660
rect 10948 16604 12460 16660
rect 12516 16604 12526 16660
rect 31714 16604 31724 16660
rect 31780 16604 33180 16660
rect 33236 16604 33246 16660
rect 11218 16492 11228 16548
rect 11284 16492 15820 16548
rect 15876 16492 15886 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 18722 16380 18732 16436
rect 18788 16380 19516 16436
rect 19572 16380 19582 16436
rect 12562 16268 12572 16324
rect 12628 16268 13468 16324
rect 13524 16268 13534 16324
rect 17490 16268 17500 16324
rect 17556 16268 18172 16324
rect 18228 16268 18620 16324
rect 18676 16268 18686 16324
rect 34626 16268 34636 16324
rect 34692 16268 39004 16324
rect 39060 16268 39070 16324
rect 0 16212 800 16240
rect 41200 16212 42000 16240
rect 0 16156 2156 16212
rect 2212 16156 2222 16212
rect 2930 16156 2940 16212
rect 2996 16156 13580 16212
rect 13636 16156 13646 16212
rect 19394 16156 19404 16212
rect 19460 16156 21084 16212
rect 21140 16156 21150 16212
rect 33282 16156 33292 16212
rect 33348 16156 35532 16212
rect 35588 16156 35598 16212
rect 39778 16156 39788 16212
rect 39844 16156 42000 16212
rect 0 16128 800 16156
rect 41200 16128 42000 16156
rect 18386 16044 18396 16100
rect 18452 16044 19292 16100
rect 19348 16044 20188 16100
rect 20244 16044 20254 16100
rect 20514 16044 20524 16100
rect 20580 16044 21308 16100
rect 21364 16044 23996 16100
rect 24052 16044 26684 16100
rect 26740 16044 28588 16100
rect 28644 16044 29260 16100
rect 29316 16044 29326 16100
rect 29586 16044 29596 16100
rect 29652 16044 30268 16100
rect 30324 16044 30334 16100
rect 31602 16044 31612 16100
rect 31668 16044 39004 16100
rect 39060 16044 39070 16100
rect 11106 15932 11116 15988
rect 11172 15932 11900 15988
rect 11956 15932 11966 15988
rect 26002 15932 26012 15988
rect 26068 15932 27244 15988
rect 27300 15932 29932 15988
rect 29988 15932 31052 15988
rect 31108 15932 31118 15988
rect 33282 15932 33292 15988
rect 33348 15932 34524 15988
rect 34580 15932 34590 15988
rect 15092 15820 21196 15876
rect 21252 15820 21262 15876
rect 26338 15820 26348 15876
rect 26404 15820 26908 15876
rect 26964 15820 26974 15876
rect 28130 15820 28140 15876
rect 28196 15820 29260 15876
rect 29316 15820 29326 15876
rect 30706 15820 30716 15876
rect 30772 15820 32396 15876
rect 32452 15820 33404 15876
rect 33460 15820 33470 15876
rect 33954 15820 33964 15876
rect 34020 15820 35084 15876
rect 35140 15820 35532 15876
rect 35588 15820 35598 15876
rect 0 15540 800 15568
rect 0 15484 2044 15540
rect 2100 15484 2110 15540
rect 9538 15484 9548 15540
rect 9604 15484 10108 15540
rect 10164 15484 10174 15540
rect 13570 15484 13580 15540
rect 13636 15484 14364 15540
rect 14420 15484 14430 15540
rect 0 15456 800 15484
rect 10108 15428 10164 15484
rect 15092 15428 15148 15820
rect 32050 15708 32060 15764
rect 32116 15708 32956 15764
rect 33012 15708 33022 15764
rect 34402 15708 34412 15764
rect 34468 15708 34860 15764
rect 34916 15708 39228 15764
rect 39284 15708 39294 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 29810 15596 29820 15652
rect 29876 15596 32284 15652
rect 32340 15596 32350 15652
rect 41200 15540 42000 15568
rect 17490 15484 17500 15540
rect 17556 15484 18396 15540
rect 18452 15484 18462 15540
rect 24658 15484 24668 15540
rect 24724 15484 25788 15540
rect 25844 15484 25854 15540
rect 32162 15484 32172 15540
rect 32228 15484 39116 15540
rect 39172 15484 39182 15540
rect 40114 15484 40124 15540
rect 40180 15484 42000 15540
rect 41200 15456 42000 15484
rect 10108 15372 14476 15428
rect 14532 15372 15148 15428
rect 19170 15372 19180 15428
rect 19236 15372 22148 15428
rect 31154 15372 31164 15428
rect 31220 15372 33740 15428
rect 33796 15372 33806 15428
rect 22092 15316 22148 15372
rect 32620 15316 32676 15372
rect 16258 15260 16268 15316
rect 16324 15260 17276 15316
rect 17332 15260 17342 15316
rect 19618 15260 19628 15316
rect 19684 15260 20860 15316
rect 20916 15260 20926 15316
rect 22082 15260 22092 15316
rect 22148 15260 23324 15316
rect 23380 15260 25340 15316
rect 25396 15260 25406 15316
rect 26898 15260 26908 15316
rect 26964 15260 31052 15316
rect 31108 15260 32060 15316
rect 32116 15260 32126 15316
rect 32610 15260 32620 15316
rect 32676 15260 32686 15316
rect 33618 15260 33628 15316
rect 33684 15260 34636 15316
rect 34692 15260 34702 15316
rect 33628 15204 33684 15260
rect 15362 15148 15372 15204
rect 15428 15148 16716 15204
rect 16772 15148 18060 15204
rect 18116 15148 18126 15204
rect 18722 15148 18732 15204
rect 18788 15148 19740 15204
rect 19796 15148 19806 15204
rect 21308 15148 25676 15204
rect 25732 15148 25742 15204
rect 30818 15148 30828 15204
rect 30884 15148 31500 15204
rect 31556 15148 31566 15204
rect 31892 15148 33684 15204
rect 17948 15092 18004 15148
rect 17948 15036 19068 15092
rect 19124 15036 19134 15092
rect 18508 14980 18564 15036
rect 21308 14980 21364 15148
rect 31892 15092 31948 15148
rect 31042 15036 31052 15092
rect 31108 15036 31948 15092
rect 33170 15036 33180 15092
rect 33236 15036 34748 15092
rect 34804 15036 35756 15092
rect 35812 15036 35822 15092
rect 18498 14924 18508 14980
rect 18564 14924 18574 14980
rect 21298 14924 21308 14980
rect 21364 14924 21374 14980
rect 32610 14924 32620 14980
rect 32676 14924 33292 14980
rect 33348 14924 34636 14980
rect 34692 14924 34702 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 41200 14868 42000 14896
rect 19058 14812 19068 14868
rect 19124 14812 26124 14868
rect 26180 14812 26190 14868
rect 30594 14812 30604 14868
rect 30660 14812 31500 14868
rect 31556 14812 31566 14868
rect 39778 14812 39788 14868
rect 39844 14812 42000 14868
rect 41200 14784 42000 14812
rect 21522 14700 21532 14756
rect 21588 14700 21868 14756
rect 21924 14700 21934 14756
rect 27122 14700 27132 14756
rect 27188 14700 27580 14756
rect 27636 14700 27646 14756
rect 27906 14700 27916 14756
rect 27972 14700 39004 14756
rect 39060 14700 39070 14756
rect 19282 14588 19292 14644
rect 19348 14588 22540 14644
rect 22596 14588 26236 14644
rect 26292 14588 26302 14644
rect 27234 14588 27244 14644
rect 27300 14588 28028 14644
rect 28084 14588 30716 14644
rect 30772 14588 30782 14644
rect 10098 14476 10108 14532
rect 10164 14476 10668 14532
rect 10724 14476 13692 14532
rect 13748 14476 14252 14532
rect 14308 14476 14924 14532
rect 14980 14476 14990 14532
rect 20178 14476 20188 14532
rect 20244 14476 22204 14532
rect 22260 14476 24780 14532
rect 24836 14476 24846 14532
rect 26114 14476 26124 14532
rect 26180 14476 27020 14532
rect 27076 14476 27086 14532
rect 29698 14476 29708 14532
rect 29764 14476 31052 14532
rect 31108 14476 31118 14532
rect 7522 14364 7532 14420
rect 7588 14364 8428 14420
rect 8484 14364 8494 14420
rect 21634 14364 21644 14420
rect 21700 14364 23212 14420
rect 23268 14364 23996 14420
rect 24052 14364 24062 14420
rect 26562 14364 26572 14420
rect 26628 14364 28252 14420
rect 28308 14364 28924 14420
rect 28980 14364 28990 14420
rect 32946 14364 32956 14420
rect 33012 14364 34188 14420
rect 34244 14364 34254 14420
rect 7186 14252 7196 14308
rect 7252 14252 7868 14308
rect 7924 14252 7934 14308
rect 27010 14252 27020 14308
rect 27076 14252 27916 14308
rect 27972 14252 27982 14308
rect 28354 14252 28364 14308
rect 28420 14252 30940 14308
rect 30996 14252 31006 14308
rect 34850 14252 34860 14308
rect 34916 14252 36092 14308
rect 36148 14252 36158 14308
rect 41200 14196 42000 14224
rect 25218 14140 25228 14196
rect 25284 14140 27356 14196
rect 27412 14140 27422 14196
rect 40226 14140 40236 14196
rect 40292 14140 42000 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 41200 14112 42000 14140
rect 15922 13916 15932 13972
rect 15988 13916 16828 13972
rect 16884 13916 22428 13972
rect 22484 13916 22494 13972
rect 24098 13916 24108 13972
rect 24164 13916 26796 13972
rect 26852 13916 26862 13972
rect 30380 13916 33068 13972
rect 33124 13916 33134 13972
rect 34178 13916 34188 13972
rect 34244 13916 38556 13972
rect 38612 13916 38622 13972
rect 2930 13804 2940 13860
rect 2996 13804 5068 13860
rect 5124 13804 5134 13860
rect 16370 13804 16380 13860
rect 16436 13804 17836 13860
rect 17892 13804 21308 13860
rect 21364 13804 21374 13860
rect 23762 13804 23772 13860
rect 23828 13804 28140 13860
rect 28196 13804 29148 13860
rect 29204 13804 29214 13860
rect 8978 13692 8988 13748
rect 9044 13692 9660 13748
rect 9716 13692 9726 13748
rect 6066 13580 6076 13636
rect 6132 13580 7196 13636
rect 7252 13580 7262 13636
rect 21410 13580 21420 13636
rect 21476 13580 23884 13636
rect 23940 13580 23950 13636
rect 24322 13580 24332 13636
rect 24388 13580 25452 13636
rect 25508 13580 25518 13636
rect 26572 13580 26908 13636
rect 27010 13580 27020 13636
rect 27076 13580 28028 13636
rect 28084 13580 28094 13636
rect 26572 13524 26628 13580
rect 18834 13468 18844 13524
rect 18900 13468 19292 13524
rect 19348 13468 19358 13524
rect 24210 13468 24220 13524
rect 24276 13468 26628 13524
rect 26852 13524 26908 13580
rect 30380 13524 30436 13916
rect 30594 13804 30604 13860
rect 30660 13804 32508 13860
rect 32564 13804 32574 13860
rect 30930 13692 30940 13748
rect 30996 13692 31612 13748
rect 31668 13692 32284 13748
rect 32340 13692 32732 13748
rect 32788 13692 35644 13748
rect 35700 13692 38668 13748
rect 38724 13692 38734 13748
rect 32050 13580 32060 13636
rect 32116 13580 32844 13636
rect 32900 13580 34524 13636
rect 34580 13580 34590 13636
rect 41200 13524 42000 13552
rect 26852 13468 30380 13524
rect 30436 13468 30446 13524
rect 31154 13468 31164 13524
rect 31220 13468 34076 13524
rect 34132 13468 34142 13524
rect 40002 13468 40012 13524
rect 40068 13468 42000 13524
rect 41200 13440 42000 13468
rect 26012 13356 27020 13412
rect 27076 13356 27086 13412
rect 27234 13356 27244 13412
rect 27300 13356 28140 13412
rect 28196 13356 29596 13412
rect 29652 13356 29662 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 26012 13188 26068 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 5058 13132 5068 13188
rect 5124 13132 6524 13188
rect 6580 13132 7308 13188
rect 7364 13132 7374 13188
rect 23492 13132 23772 13188
rect 23828 13132 23838 13188
rect 26002 13132 26012 13188
rect 26068 13132 26078 13188
rect 26226 13132 26236 13188
rect 26292 13132 26908 13188
rect 26964 13132 26974 13188
rect 28018 13132 28028 13188
rect 28084 13132 29708 13188
rect 29764 13132 29774 13188
rect 30482 13132 30492 13188
rect 30548 13132 30828 13188
rect 30884 13132 30894 13188
rect 32722 13132 32732 13188
rect 32788 13132 33516 13188
rect 33572 13132 33582 13188
rect 34178 13132 34188 13188
rect 34244 13132 35532 13188
rect 35588 13132 35598 13188
rect 23492 13076 23548 13132
rect 10882 13020 10892 13076
rect 10948 13020 12012 13076
rect 12068 13020 12078 13076
rect 14690 13020 14700 13076
rect 14756 13020 15260 13076
rect 15316 13020 15326 13076
rect 15586 13020 15596 13076
rect 15652 13020 18508 13076
rect 18564 13020 18574 13076
rect 20402 13020 20412 13076
rect 20468 13020 23548 13076
rect 24770 13020 24780 13076
rect 24836 13020 25676 13076
rect 25732 13020 25742 13076
rect 25900 13020 27132 13076
rect 27188 13020 27198 13076
rect 27458 13020 27468 13076
rect 27524 13020 30716 13076
rect 30772 13020 30782 13076
rect 2258 12908 2268 12964
rect 2324 12908 4844 12964
rect 4900 12908 7980 12964
rect 8036 12908 8540 12964
rect 8596 12908 8606 12964
rect 20514 12908 20524 12964
rect 20580 12908 21084 12964
rect 21140 12908 22092 12964
rect 22148 12908 22158 12964
rect 22866 12908 22876 12964
rect 22932 12908 25340 12964
rect 25396 12908 25406 12964
rect 25900 12852 25956 13020
rect 28476 12964 28532 13020
rect 26338 12908 26348 12964
rect 26404 12908 27804 12964
rect 27860 12908 27870 12964
rect 28354 12908 28364 12964
rect 28420 12908 28532 12964
rect 34738 12908 34748 12964
rect 34804 12908 35980 12964
rect 36036 12908 36046 12964
rect 41200 12852 42000 12880
rect 7634 12796 7644 12852
rect 7700 12796 8764 12852
rect 8820 12796 8830 12852
rect 18498 12796 18508 12852
rect 18564 12796 21868 12852
rect 21924 12796 22652 12852
rect 22708 12796 25228 12852
rect 25284 12796 25294 12852
rect 25442 12796 25452 12852
rect 25508 12796 25956 12852
rect 27570 12796 27580 12852
rect 27636 12796 33068 12852
rect 33124 12796 33134 12852
rect 34514 12796 34524 12852
rect 34580 12796 34972 12852
rect 35028 12796 35038 12852
rect 39442 12796 39452 12852
rect 39508 12796 40236 12852
rect 40292 12796 42000 12852
rect 41200 12768 42000 12796
rect 11218 12684 11228 12740
rect 11284 12684 11900 12740
rect 11956 12684 11966 12740
rect 26002 12684 26012 12740
rect 26068 12684 26684 12740
rect 26740 12684 26750 12740
rect 27122 12684 27132 12740
rect 27188 12684 28140 12740
rect 28196 12684 28206 12740
rect 34178 12684 34188 12740
rect 34244 12684 34636 12740
rect 34692 12684 36204 12740
rect 36260 12684 36270 12740
rect 28018 12572 28028 12628
rect 28084 12572 28812 12628
rect 28868 12572 28878 12628
rect 29362 12572 29372 12628
rect 29428 12572 30604 12628
rect 30660 12572 30670 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 33618 12348 33628 12404
rect 33684 12348 34524 12404
rect 34580 12348 34590 12404
rect 35970 12348 35980 12404
rect 36036 12348 39676 12404
rect 39732 12348 39742 12404
rect 8530 12236 8540 12292
rect 8596 12236 9996 12292
rect 10052 12236 10062 12292
rect 20290 12236 20300 12292
rect 20356 12236 22988 12292
rect 23044 12236 23772 12292
rect 23828 12236 23838 12292
rect 28914 12236 28924 12292
rect 28980 12236 29932 12292
rect 29988 12236 29998 12292
rect 30594 12236 30604 12292
rect 30660 12236 33740 12292
rect 33796 12236 33806 12292
rect 34066 12236 34076 12292
rect 34132 12236 34972 12292
rect 35028 12236 35038 12292
rect 33740 12180 33796 12236
rect 20850 12124 20860 12180
rect 20916 12124 22204 12180
rect 22260 12124 22270 12180
rect 25218 12124 25228 12180
rect 25284 12124 25452 12180
rect 25508 12124 25518 12180
rect 28466 12124 28476 12180
rect 28532 12124 29596 12180
rect 29652 12124 29662 12180
rect 30034 12124 30044 12180
rect 30100 12124 30716 12180
rect 30772 12124 30782 12180
rect 33740 12124 34748 12180
rect 34804 12124 34814 12180
rect 22754 12012 22764 12068
rect 22820 12012 24556 12068
rect 24612 12012 24622 12068
rect 26674 12012 26684 12068
rect 26740 12012 27020 12068
rect 27076 12012 27086 12068
rect 30818 12012 30828 12068
rect 30884 12012 34636 12068
rect 34692 12012 34702 12068
rect 11330 11900 11340 11956
rect 11396 11900 13580 11956
rect 13636 11900 13646 11956
rect 19954 11900 19964 11956
rect 20020 11900 22876 11956
rect 22932 11900 23660 11956
rect 23716 11900 23726 11956
rect 26450 11900 26460 11956
rect 26516 11900 27244 11956
rect 27300 11900 27310 11956
rect 32050 11900 32060 11956
rect 32116 11900 33964 11956
rect 34020 11900 35196 11956
rect 35252 11900 35532 11956
rect 35588 11900 35980 11956
rect 36036 11900 36046 11956
rect 19842 11788 19852 11844
rect 19908 11788 20412 11844
rect 20468 11788 23100 11844
rect 23156 11788 23166 11844
rect 31892 11788 34076 11844
rect 34132 11788 34142 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 31892 11732 31948 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 16706 11676 16716 11732
rect 16772 11676 19628 11732
rect 19684 11676 19694 11732
rect 28242 11676 28252 11732
rect 28308 11676 29484 11732
rect 29540 11676 31948 11732
rect 5954 11564 5964 11620
rect 6020 11564 6860 11620
rect 6916 11564 6926 11620
rect 12898 11452 12908 11508
rect 12964 11452 14364 11508
rect 14420 11452 14430 11508
rect 18050 11452 18060 11508
rect 18116 11452 18732 11508
rect 18788 11452 18798 11508
rect 26898 11452 26908 11508
rect 26964 11452 27692 11508
rect 27748 11452 27758 11508
rect 30930 11452 30940 11508
rect 30996 11452 33404 11508
rect 33460 11452 33470 11508
rect 28466 11340 28476 11396
rect 28532 11340 29820 11396
rect 29876 11340 30380 11396
rect 30436 11340 30446 11396
rect 31154 11340 31164 11396
rect 31220 11340 31836 11396
rect 31892 11340 31902 11396
rect 33730 11340 33740 11396
rect 33796 11340 34524 11396
rect 34580 11340 34972 11396
rect 35028 11340 36148 11396
rect 36092 11284 36148 11340
rect 10770 11228 10780 11284
rect 10836 11228 13916 11284
rect 13972 11228 13982 11284
rect 20962 11228 20972 11284
rect 21028 11228 21868 11284
rect 21924 11228 21934 11284
rect 24434 11228 24444 11284
rect 24500 11228 25228 11284
rect 25284 11228 25294 11284
rect 30594 11228 30604 11284
rect 30660 11228 31052 11284
rect 31108 11228 31118 11284
rect 31266 11228 31276 11284
rect 31332 11228 31342 11284
rect 33954 11228 33964 11284
rect 34020 11228 35084 11284
rect 35140 11228 35150 11284
rect 36082 11228 36092 11284
rect 36148 11228 37212 11284
rect 37268 11228 37278 11284
rect 31276 11172 31332 11228
rect 9650 11116 9660 11172
rect 9716 11116 10332 11172
rect 10388 11116 10398 11172
rect 28242 11116 28252 11172
rect 28308 11116 29260 11172
rect 29316 11116 29326 11172
rect 31276 11116 34300 11172
rect 34356 11116 34366 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 30930 10780 30940 10836
rect 30996 10780 31276 10836
rect 31332 10780 31342 10836
rect 23762 10668 23772 10724
rect 23828 10668 25340 10724
rect 25396 10668 25406 10724
rect 28354 10668 28364 10724
rect 28420 10668 31612 10724
rect 31668 10668 31678 10724
rect 37650 10668 37660 10724
rect 37716 10668 38668 10724
rect 38724 10668 39116 10724
rect 39172 10668 39182 10724
rect 11442 10444 11452 10500
rect 11508 10444 12460 10500
rect 12516 10444 12526 10500
rect 22194 10444 22204 10500
rect 22260 10444 22876 10500
rect 22932 10444 22942 10500
rect 24994 10332 25004 10388
rect 25060 10332 25900 10388
rect 25956 10332 30604 10388
rect 30660 10332 32284 10388
rect 32340 10332 34300 10388
rect 34356 10332 35308 10388
rect 35364 10332 35374 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 9426 9996 9436 10052
rect 9492 9996 10780 10052
rect 10836 9996 10846 10052
rect 19730 9996 19740 10052
rect 19796 9996 20972 10052
rect 21028 9996 21038 10052
rect 25106 9996 25116 10052
rect 25172 9996 27132 10052
rect 27188 9996 27198 10052
rect 27570 9996 27580 10052
rect 27636 9996 30044 10052
rect 30100 9996 30110 10052
rect 32050 9996 32060 10052
rect 32116 9996 34636 10052
rect 34692 9996 34702 10052
rect 30044 9940 30100 9996
rect 12562 9884 12572 9940
rect 12628 9884 13020 9940
rect 13076 9884 13692 9940
rect 13748 9884 15372 9940
rect 15428 9884 15438 9940
rect 18834 9884 18844 9940
rect 18900 9884 21644 9940
rect 21700 9884 21710 9940
rect 24770 9884 24780 9940
rect 24836 9884 26460 9940
rect 26516 9884 26526 9940
rect 30044 9884 33516 9940
rect 33572 9884 33582 9940
rect 20738 9772 20748 9828
rect 20804 9772 21308 9828
rect 21364 9772 21868 9828
rect 21924 9772 21934 9828
rect 24322 9772 24332 9828
rect 24388 9772 25452 9828
rect 25508 9772 25518 9828
rect 26562 9772 26572 9828
rect 26628 9772 27020 9828
rect 27076 9772 27086 9828
rect 29250 9772 29260 9828
rect 29316 9772 30156 9828
rect 30212 9772 30222 9828
rect 33954 9772 33964 9828
rect 34020 9772 35532 9828
rect 35588 9772 35598 9828
rect 20514 9660 20524 9716
rect 20580 9660 22428 9716
rect 22484 9660 22494 9716
rect 23202 9660 23212 9716
rect 23268 9660 30716 9716
rect 30772 9660 30782 9716
rect 31490 9660 31500 9716
rect 31556 9660 32284 9716
rect 32340 9660 32350 9716
rect 32834 9660 32844 9716
rect 32900 9660 34188 9716
rect 34244 9660 34636 9716
rect 34692 9660 36316 9716
rect 36372 9660 36382 9716
rect 32844 9604 32900 9660
rect 19618 9548 19628 9604
rect 19684 9548 21420 9604
rect 21476 9548 21486 9604
rect 25218 9548 25228 9604
rect 25284 9548 26796 9604
rect 26852 9548 26862 9604
rect 30034 9548 30044 9604
rect 30100 9548 30828 9604
rect 30884 9548 30894 9604
rect 31938 9548 31948 9604
rect 32004 9548 32900 9604
rect 34738 9548 34748 9604
rect 34804 9548 36204 9604
rect 36260 9548 36270 9604
rect 27122 9436 27132 9492
rect 27188 9436 29372 9492
rect 29428 9436 29438 9492
rect 30930 9436 30940 9492
rect 30996 9436 31388 9492
rect 31444 9436 31454 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 34748 9380 34804 9548
rect 25890 9324 25900 9380
rect 25956 9324 29260 9380
rect 29316 9324 29326 9380
rect 29586 9324 29596 9380
rect 29652 9324 34804 9380
rect 24770 9212 24780 9268
rect 24836 9212 26012 9268
rect 26068 9212 26078 9268
rect 28914 9212 28924 9268
rect 28980 9212 30380 9268
rect 30436 9212 30446 9268
rect 32274 9212 32284 9268
rect 32340 9212 34076 9268
rect 34132 9212 35084 9268
rect 35140 9212 35150 9268
rect 26450 9100 26460 9156
rect 26516 9100 26908 9156
rect 26964 9100 28476 9156
rect 28532 9100 29372 9156
rect 29428 9100 29438 9156
rect 31490 9100 31500 9156
rect 31556 9100 33852 9156
rect 33908 9100 33918 9156
rect 31602 8988 31612 9044
rect 31668 8988 32060 9044
rect 32116 8988 32126 9044
rect 32610 8988 32620 9044
rect 32676 8988 33964 9044
rect 34020 8988 34030 9044
rect 31826 8876 31836 8932
rect 31892 8876 33068 8932
rect 33124 8876 33134 8932
rect 29698 8764 29708 8820
rect 29764 8764 30268 8820
rect 30324 8764 31500 8820
rect 31556 8764 31566 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 29362 8316 29372 8372
rect 29428 8316 30604 8372
rect 30660 8316 30940 8372
rect 30996 8316 31006 8372
rect 31154 8316 31164 8372
rect 31220 8316 31724 8372
rect 31780 8316 31790 8372
rect 28130 8204 28140 8260
rect 28196 8204 29148 8260
rect 29204 8204 29214 8260
rect 31266 8204 31276 8260
rect 31332 8204 32620 8260
rect 32676 8204 33068 8260
rect 33124 8204 33134 8260
rect 27458 8092 27468 8148
rect 27524 8092 28028 8148
rect 28084 8092 31948 8148
rect 32004 8092 32014 8148
rect 25106 7980 25116 8036
rect 25172 7980 25900 8036
rect 25956 7980 25966 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 22642 7532 22652 7588
rect 22708 7532 23436 7588
rect 23492 7532 23502 7588
rect 23762 7532 23772 7588
rect 23828 7532 25340 7588
rect 25396 7532 25406 7588
rect 28690 7532 28700 7588
rect 28756 7532 31836 7588
rect 31892 7532 31902 7588
rect 32386 7532 32396 7588
rect 32452 7532 35420 7588
rect 35476 7532 35868 7588
rect 35924 7532 37660 7588
rect 37716 7532 37726 7588
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 22194 6636 22204 6692
rect 22260 6636 23772 6692
rect 23828 6636 25788 6692
rect 25844 6636 28364 6692
rect 28420 6636 31724 6692
rect 31780 6636 31790 6692
rect 26786 6524 26796 6580
rect 26852 6524 27804 6580
rect 27860 6524 27870 6580
rect 22418 6412 22428 6468
rect 22484 6412 26012 6468
rect 26068 6412 27916 6468
rect 27972 6412 27982 6468
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 18162 3612 18172 3668
rect 18228 3612 18844 3668
rect 18900 3612 18910 3668
rect 23090 3500 23100 3556
rect 23156 3500 23548 3556
rect 23604 3500 23614 3556
rect 21074 3388 21084 3444
rect 21140 3388 21756 3444
rect 21812 3388 21822 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0595_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21280 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0596_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23296 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0597_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19824 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0598_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19936 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0599_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0600_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18144 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0601_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _0602_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20160 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _0603_
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0604_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21280 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0605_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0606_
timestamp 1698431365
transform -1 0 17808 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0607_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15120 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0608_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0609_
timestamp 1698431365
transform -1 0 17808 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0610_
timestamp 1698431365
transform 1 0 15456 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0611_
timestamp 1698431365
transform -1 0 23520 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0612_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22176 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0613_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0614_
timestamp 1698431365
transform 1 0 26656 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0615_
timestamp 1698431365
transform -1 0 27440 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0616_
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _0617_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0618_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0619_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23968 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0620_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30912 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0621_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0622_
timestamp 1698431365
transform -1 0 28336 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0623_
timestamp 1698431365
transform -1 0 34832 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0624_
timestamp 1698431365
transform 1 0 33824 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0625_
timestamp 1698431365
transform 1 0 33488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0626_
timestamp 1698431365
transform 1 0 32480 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0627_
timestamp 1698431365
transform -1 0 33488 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0628_
timestamp 1698431365
transform 1 0 30912 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0629_
timestamp 1698431365
transform -1 0 19040 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_4  _0630_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18480 0 1 15680
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0631_
timestamp 1698431365
transform 1 0 31360 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0632_
timestamp 1698431365
transform -1 0 33488 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0633_
timestamp 1698431365
transform 1 0 19152 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0634_
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0635_
timestamp 1698431365
transform -1 0 18144 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0636_
timestamp 1698431365
transform 1 0 17360 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0637_
timestamp 1698431365
transform 1 0 16016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0638_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16240 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0639_
timestamp 1698431365
transform -1 0 18592 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0640_
timestamp 1698431365
transform -1 0 14896 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0641_
timestamp 1698431365
transform -1 0 14224 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0642_
timestamp 1698431365
transform 1 0 8512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0643_
timestamp 1698431365
transform 1 0 9296 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _0644_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12544 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0645_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12432 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0646_
timestamp 1698431365
transform 1 0 7840 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0647_
timestamp 1698431365
transform -1 0 12208 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0648_
timestamp 1698431365
transform 1 0 11312 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0649_
timestamp 1698431365
transform 1 0 7168 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0650_
timestamp 1698431365
transform 1 0 9072 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0651_
timestamp 1698431365
transform 1 0 8512 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0652_
timestamp 1698431365
transform 1 0 8624 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0653_
timestamp 1698431365
transform 1 0 8400 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0654_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8624 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0655_
timestamp 1698431365
transform -1 0 13888 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0656_
timestamp 1698431365
transform -1 0 14336 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _0657_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11872 0 -1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0658_
timestamp 1698431365
transform -1 0 15680 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0659_
timestamp 1698431365
transform -1 0 19936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0660_
timestamp 1698431365
transform -1 0 16128 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0661_
timestamp 1698431365
transform -1 0 19152 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0662_
timestamp 1698431365
transform -1 0 15120 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0663_
timestamp 1698431365
transform 1 0 14560 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0664_
timestamp 1698431365
transform -1 0 18480 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0665_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18368 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0666_
timestamp 1698431365
transform 1 0 20496 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _0667_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12880 0 1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0668_
timestamp 1698431365
transform 1 0 7392 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0669_
timestamp 1698431365
transform 1 0 6944 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _0670_
timestamp 1698431365
transform 1 0 6048 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _0671_
timestamp 1698431365
transform 1 0 5936 0 -1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0672_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0673_
timestamp 1698431365
transform -1 0 11312 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0674_
timestamp 1698431365
transform -1 0 13888 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0675_
timestamp 1698431365
transform 1 0 10304 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0676_
timestamp 1698431365
transform 1 0 11648 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0677_
timestamp 1698431365
transform -1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0678_
timestamp 1698431365
transform 1 0 14224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0679_
timestamp 1698431365
transform 1 0 15680 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0680_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17360 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0681_
timestamp 1698431365
transform 1 0 14784 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0682_
timestamp 1698431365
transform -1 0 12768 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0683_
timestamp 1698431365
transform -1 0 13776 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0684_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11648 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0685_
timestamp 1698431365
transform -1 0 12544 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0686_
timestamp 1698431365
transform 1 0 11536 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0687_
timestamp 1698431365
transform -1 0 25760 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0688_
timestamp 1698431365
transform 1 0 22176 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0689_
timestamp 1698431365
transform 1 0 19824 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0690_
timestamp 1698431365
transform 1 0 19600 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0691_
timestamp 1698431365
transform 1 0 24192 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _0692_
timestamp 1698431365
transform -1 0 26432 0 1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0693_
timestamp 1698431365
transform -1 0 30912 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0694_
timestamp 1698431365
transform 1 0 27664 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0695_
timestamp 1698431365
transform -1 0 35952 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _0696_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29792 0 1 23520
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0697_
timestamp 1698431365
transform -1 0 34720 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0698_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33152 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0699_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34944 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0700_
timestamp 1698431365
transform -1 0 34944 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0701_
timestamp 1698431365
transform 1 0 30464 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0702_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0703_
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0704_
timestamp 1698431365
transform -1 0 30464 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0705_
timestamp 1698431365
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _0706_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32368 0 -1 23520
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0707_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0708_
timestamp 1698431365
transform -1 0 26432 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0709_
timestamp 1698431365
transform -1 0 24528 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0710_
timestamp 1698431365
transform -1 0 27888 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0711_
timestamp 1698431365
transform 1 0 25200 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0712_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27776 0 -1 21952
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0713_
timestamp 1698431365
transform -1 0 24192 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0714_
timestamp 1698431365
transform 1 0 20048 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0715_
timestamp 1698431365
transform 1 0 22848 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0716_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22176 0 1 23520
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _0717_
timestamp 1698431365
transform -1 0 26768 0 1 21952
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0718_
timestamp 1698431365
transform 1 0 14784 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0719_
timestamp 1698431365
transform -1 0 17024 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0720_
timestamp 1698431365
transform -1 0 15680 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0721_
timestamp 1698431365
transform 1 0 11984 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0722_
timestamp 1698431365
transform -1 0 11648 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0723_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14000 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0724_
timestamp 1698431365
transform 1 0 9744 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0725_
timestamp 1698431365
transform -1 0 6496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0726_
timestamp 1698431365
transform -1 0 6048 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0727_
timestamp 1698431365
transform 1 0 6048 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0728_
timestamp 1698431365
transform -1 0 6720 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0729_
timestamp 1698431365
transform 1 0 6720 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0730_
timestamp 1698431365
transform 1 0 6048 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0731_
timestamp 1698431365
transform 1 0 9744 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0732_
timestamp 1698431365
transform 1 0 12432 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0733_
timestamp 1698431365
transform 1 0 8512 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0734_
timestamp 1698431365
transform 1 0 10976 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0735_
timestamp 1698431365
transform 1 0 11088 0 -1 25088
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0736_
timestamp 1698431365
transform 1 0 7280 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0737_
timestamp 1698431365
transform 1 0 7168 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0738_
timestamp 1698431365
transform -1 0 11200 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0739_
timestamp 1698431365
transform -1 0 10752 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0740_
timestamp 1698431365
transform 1 0 11760 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0741_
timestamp 1698431365
transform -1 0 19824 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0742_
timestamp 1698431365
transform -1 0 16688 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0743_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13664 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0744_
timestamp 1698431365
transform -1 0 14896 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0745_
timestamp 1698431365
transform 1 0 26320 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0746_
timestamp 1698431365
transform -1 0 29456 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0747_
timestamp 1698431365
transform 1 0 25984 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0748_
timestamp 1698431365
transform -1 0 29120 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0749_
timestamp 1698431365
transform -1 0 26208 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0750_
timestamp 1698431365
transform -1 0 24864 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0751_
timestamp 1698431365
transform 1 0 22624 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0752_
timestamp 1698431365
transform 1 0 21504 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0753_
timestamp 1698431365
transform 1 0 22512 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0754_
timestamp 1698431365
transform 1 0 23072 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0755_
timestamp 1698431365
transform 1 0 23968 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0756_
timestamp 1698431365
transform 1 0 23072 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0757_
timestamp 1698431365
transform 1 0 25872 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0758_
timestamp 1698431365
transform -1 0 28224 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0759_
timestamp 1698431365
transform -1 0 28448 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0760_
timestamp 1698431365
transform 1 0 25984 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0761_
timestamp 1698431365
transform 1 0 23408 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0762_
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0763_
timestamp 1698431365
transform 1 0 22512 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0764_
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0765_
timestamp 1698431365
transform -1 0 25312 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0766_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26208 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0767_
timestamp 1698431365
transform -1 0 28336 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0768_
timestamp 1698431365
transform -1 0 33600 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0769_
timestamp 1698431365
transform -1 0 33488 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0770_
timestamp 1698431365
transform 1 0 33264 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0771_
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0772_
timestamp 1698431365
transform 1 0 30240 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0773_
timestamp 1698431365
transform -1 0 32032 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0774_
timestamp 1698431365
transform -1 0 34384 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0775_
timestamp 1698431365
transform 1 0 34832 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0776_
timestamp 1698431365
transform -1 0 33824 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0777_
timestamp 1698431365
transform 1 0 33600 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0778_
timestamp 1698431365
transform -1 0 35952 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0779_
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0780_
timestamp 1698431365
transform -1 0 32704 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0781_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0782_
timestamp 1698431365
transform -1 0 31360 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0783_
timestamp 1698431365
transform 1 0 17920 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0784_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0785_
timestamp 1698431365
transform 1 0 21840 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0786_
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0787_
timestamp 1698431365
transform 1 0 7952 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _0788_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30576 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0789_
timestamp 1698431365
transform -1 0 25984 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _0790_
timestamp 1698431365
transform -1 0 23520 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0791_
timestamp 1698431365
transform 1 0 12880 0 -1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0792_
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0793_
timestamp 1698431365
transform 1 0 9072 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0794_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10752 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _0795_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0796_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0797_
timestamp 1698431365
transform -1 0 17024 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0798_
timestamp 1698431365
transform 1 0 17584 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0799_
timestamp 1698431365
transform 1 0 22848 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0800_
timestamp 1698431365
transform 1 0 27776 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0801_
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0802_
timestamp 1698431365
transform 1 0 31696 0 1 29792
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0803_
timestamp 1698431365
transform -1 0 34272 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _0804_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30912 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0805_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21840 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0806_
timestamp 1698431365
transform 1 0 20160 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0807_
timestamp 1698431365
transform -1 0 20720 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0808_
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0809_
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0810_
timestamp 1698431365
transform -1 0 28336 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0811_
timestamp 1698431365
transform 1 0 30464 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0812_
timestamp 1698431365
transform 1 0 32032 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0813_
timestamp 1698431365
transform 1 0 32256 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0814_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31808 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _0815_
timestamp 1698431365
transform -1 0 35616 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0816_
timestamp 1698431365
transform -1 0 34608 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0817_
timestamp 1698431365
transform -1 0 36624 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _0818_
timestamp 1698431365
transform 1 0 19376 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0819_
timestamp 1698431365
transform -1 0 18816 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0820_
timestamp 1698431365
transform 1 0 22960 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0821_
timestamp 1698431365
transform -1 0 32256 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0822_
timestamp 1698431365
transform 1 0 30352 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0823_
timestamp 1698431365
transform 1 0 32256 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0824_
timestamp 1698431365
transform -1 0 32704 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0825_
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0826_
timestamp 1698431365
transform 1 0 30240 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0827_
timestamp 1698431365
transform 1 0 26096 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0828_
timestamp 1698431365
transform -1 0 31696 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0829_
timestamp 1698431365
transform 1 0 30464 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0830_
timestamp 1698431365
transform 1 0 26544 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0831_
timestamp 1698431365
transform -1 0 34832 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0832_
timestamp 1698431365
transform 1 0 30800 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0833_
timestamp 1698431365
transform 1 0 31248 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0834_
timestamp 1698431365
transform -1 0 33488 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0835_
timestamp 1698431365
transform 1 0 31696 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0836_
timestamp 1698431365
transform -1 0 29008 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0837_
timestamp 1698431365
transform -1 0 23072 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0838_
timestamp 1698431365
transform 1 0 23856 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0839_
timestamp 1698431365
transform 1 0 26768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0840_
timestamp 1698431365
transform -1 0 28560 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0841_
timestamp 1698431365
transform 1 0 27216 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0842_
timestamp 1698431365
transform 1 0 25536 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0843_
timestamp 1698431365
transform -1 0 24864 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0844_
timestamp 1698431365
transform 1 0 26432 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0845_
timestamp 1698431365
transform 1 0 26432 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0846_
timestamp 1698431365
transform 1 0 26768 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0847_
timestamp 1698431365
transform -1 0 28784 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0848_
timestamp 1698431365
transform 1 0 27328 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0849_
timestamp 1698431365
transform 1 0 21616 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0850_
timestamp 1698431365
transform 1 0 23856 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0851_
timestamp 1698431365
transform 1 0 23968 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0852_
timestamp 1698431365
transform 1 0 22512 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0853_
timestamp 1698431365
transform 1 0 23968 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0854_
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0855_
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0856_
timestamp 1698431365
transform 1 0 19936 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0857_
timestamp 1698431365
transform -1 0 22624 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0858_
timestamp 1698431365
transform -1 0 21952 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0859_
timestamp 1698431365
transform -1 0 22512 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0860_
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0861_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18816 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0862_
timestamp 1698431365
transform -1 0 19040 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0863_
timestamp 1698431365
transform 1 0 19600 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0864_
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0865_
timestamp 1698431365
transform 1 0 14448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0866_
timestamp 1698431365
transform 1 0 11312 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0867_
timestamp 1698431365
transform 1 0 12320 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0868_
timestamp 1698431365
transform -1 0 17808 0 1 31360
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0869_
timestamp 1698431365
transform -1 0 15792 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0870_
timestamp 1698431365
transform 1 0 17472 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0871_
timestamp 1698431365
transform 1 0 17920 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0872_
timestamp 1698431365
transform 1 0 19824 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0873_
timestamp 1698431365
transform -1 0 20272 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0874_
timestamp 1698431365
transform 1 0 20160 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0875_
timestamp 1698431365
transform 1 0 19264 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0876_
timestamp 1698431365
transform 1 0 16352 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0877_
timestamp 1698431365
transform 1 0 15008 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0878_
timestamp 1698431365
transform 1 0 16576 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0879_
timestamp 1698431365
transform 1 0 14896 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0880_
timestamp 1698431365
transform -1 0 14560 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0881_
timestamp 1698431365
transform -1 0 14336 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0882_
timestamp 1698431365
transform 1 0 14784 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0883_
timestamp 1698431365
transform 1 0 15120 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0884_
timestamp 1698431365
transform 1 0 16464 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0885_
timestamp 1698431365
transform 1 0 18368 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0886_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18816 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0887_
timestamp 1698431365
transform 1 0 16240 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0888_
timestamp 1698431365
transform 1 0 14336 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0889_
timestamp 1698431365
transform -1 0 14000 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0890_
timestamp 1698431365
transform -1 0 18032 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0891_
timestamp 1698431365
transform 1 0 14224 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0892_
timestamp 1698431365
transform 1 0 14336 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0893_
timestamp 1698431365
transform 1 0 15680 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0894_
timestamp 1698431365
transform -1 0 18592 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0895_
timestamp 1698431365
transform 1 0 16128 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0896_
timestamp 1698431365
transform 1 0 22736 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0897_
timestamp 1698431365
transform -1 0 12544 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0898_
timestamp 1698431365
transform 1 0 10864 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0899_
timestamp 1698431365
transform -1 0 11312 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0900_
timestamp 1698431365
transform 1 0 8960 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0901_
timestamp 1698431365
transform -1 0 11200 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0902_
timestamp 1698431365
transform 1 0 9856 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0903_
timestamp 1698431365
transform -1 0 12544 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0904_
timestamp 1698431365
transform 1 0 11088 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0905_
timestamp 1698431365
transform -1 0 18704 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0906_
timestamp 1698431365
transform -1 0 9072 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0907_
timestamp 1698431365
transform -1 0 8288 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0908_
timestamp 1698431365
transform 1 0 7504 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0909_
timestamp 1698431365
transform -1 0 11200 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0910_
timestamp 1698431365
transform 1 0 9744 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0911_
timestamp 1698431365
transform 1 0 8400 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0912_
timestamp 1698431365
transform -1 0 7280 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0913_
timestamp 1698431365
transform 1 0 5936 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0914_
timestamp 1698431365
transform -1 0 8400 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0915_
timestamp 1698431365
transform 1 0 9632 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0916_
timestamp 1698431365
transform -1 0 10752 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0917_
timestamp 1698431365
transform -1 0 8624 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0918_
timestamp 1698431365
transform 1 0 6160 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0919_
timestamp 1698431365
transform -1 0 6832 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0920_
timestamp 1698431365
transform 1 0 5488 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0921_
timestamp 1698431365
transform 1 0 9856 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0922_
timestamp 1698431365
transform 1 0 8512 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0923_
timestamp 1698431365
transform 1 0 9968 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0924_
timestamp 1698431365
transform -1 0 7168 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0925_
timestamp 1698431365
transform 1 0 5712 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0926_
timestamp 1698431365
transform 1 0 11648 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _0927_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 -1 23520
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0928_
timestamp 1698431365
transform 1 0 8400 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0929_
timestamp 1698431365
transform 1 0 9296 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0930_
timestamp 1698431365
transform 1 0 9968 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0931_
timestamp 1698431365
transform 1 0 9520 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0932_
timestamp 1698431365
transform 1 0 9856 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0933_
timestamp 1698431365
transform 1 0 10304 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0934_
timestamp 1698431365
transform 1 0 11424 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0935_
timestamp 1698431365
transform -1 0 13888 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0936_
timestamp 1698431365
transform 1 0 11984 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0937_
timestamp 1698431365
transform -1 0 9184 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0938_
timestamp 1698431365
transform -1 0 8512 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0939_
timestamp 1698431365
transform 1 0 7392 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0940_
timestamp 1698431365
transform -1 0 6944 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0941_
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0942_
timestamp 1698431365
transform -1 0 10640 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0943_
timestamp 1698431365
transform -1 0 7840 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0944_
timestamp 1698431365
transform 1 0 8176 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0945_
timestamp 1698431365
transform -1 0 8512 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0946_
timestamp 1698431365
transform -1 0 7728 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0947_
timestamp 1698431365
transform 1 0 6720 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0948_
timestamp 1698431365
transform 1 0 8064 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0949_
timestamp 1698431365
transform -1 0 6048 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0950_
timestamp 1698431365
transform 1 0 4368 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0951_
timestamp 1698431365
transform -1 0 9184 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0952_
timestamp 1698431365
transform -1 0 9744 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0953_
timestamp 1698431365
transform 1 0 8512 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0954_
timestamp 1698431365
transform -1 0 8960 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0955_
timestamp 1698431365
transform -1 0 5936 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0956_
timestamp 1698431365
transform 1 0 4368 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0957_
timestamp 1698431365
transform -1 0 10752 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0958_
timestamp 1698431365
transform -1 0 12992 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0959_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0960_
timestamp 1698431365
transform -1 0 14000 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0961_
timestamp 1698431365
transform -1 0 11648 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0962_
timestamp 1698431365
transform -1 0 11536 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0963_
timestamp 1698431365
transform 1 0 8176 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0964_
timestamp 1698431365
transform -1 0 10304 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0965_
timestamp 1698431365
transform 1 0 8736 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0966_
timestamp 1698431365
transform 1 0 13552 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0967_
timestamp 1698431365
transform -1 0 14448 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0968_
timestamp 1698431365
transform -1 0 13104 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0969_
timestamp 1698431365
transform 1 0 14000 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0970_
timestamp 1698431365
transform 1 0 12768 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0971_
timestamp 1698431365
transform -1 0 14448 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0972_
timestamp 1698431365
transform 1 0 11648 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0973_
timestamp 1698431365
transform -1 0 19040 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0974_
timestamp 1698431365
transform 1 0 16016 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0975_
timestamp 1698431365
transform 1 0 18480 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0976_
timestamp 1698431365
transform 1 0 16016 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0977_
timestamp 1698431365
transform 1 0 17920 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0978_
timestamp 1698431365
transform 1 0 14672 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0979_
timestamp 1698431365
transform -1 0 18256 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0980_
timestamp 1698431365
transform -1 0 18368 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0981_
timestamp 1698431365
transform -1 0 17136 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0982_
timestamp 1698431365
transform 1 0 14224 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0983_
timestamp 1698431365
transform -1 0 17920 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0984_
timestamp 1698431365
transform 1 0 15456 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0985_
timestamp 1698431365
transform 1 0 16800 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0986_
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0987_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0988_
timestamp 1698431365
transform -1 0 24416 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0989_
timestamp 1698431365
transform -1 0 22624 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0990_
timestamp 1698431365
transform 1 0 21504 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0991_
timestamp 1698431365
transform -1 0 26432 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0992_
timestamp 1698431365
transform -1 0 21504 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0993_
timestamp 1698431365
transform 1 0 21280 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0994_
timestamp 1698431365
transform 1 0 21280 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0995_
timestamp 1698431365
transform -1 0 23632 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0996_
timestamp 1698431365
transform -1 0 24080 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0997_
timestamp 1698431365
transform 1 0 22624 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0998_
timestamp 1698431365
transform -1 0 20944 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0999_
timestamp 1698431365
transform -1 0 21952 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1000_
timestamp 1698431365
transform -1 0 22288 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1001_
timestamp 1698431365
transform 1 0 20272 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1002_
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1003_
timestamp 1698431365
transform -1 0 19936 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1004_
timestamp 1698431365
transform 1 0 18480 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1005_
timestamp 1698431365
transform -1 0 26992 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1006_
timestamp 1698431365
transform 1 0 23520 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1007_
timestamp 1698431365
transform 1 0 26432 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1008_
timestamp 1698431365
transform -1 0 24864 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1009_
timestamp 1698431365
transform 1 0 25984 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1010_
timestamp 1698431365
transform 1 0 23520 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1011_
timestamp 1698431365
transform -1 0 21952 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1012_
timestamp 1698431365
transform -1 0 30352 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1013_
timestamp 1698431365
transform -1 0 28112 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1014_
timestamp 1698431365
transform -1 0 29120 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1015_
timestamp 1698431365
transform 1 0 26656 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1016_
timestamp 1698431365
transform 1 0 25648 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1017_
timestamp 1698431365
transform -1 0 27104 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1018_
timestamp 1698431365
transform 1 0 34384 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1019_
timestamp 1698431365
transform -1 0 36512 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1020_
timestamp 1698431365
transform 1 0 31920 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1021_
timestamp 1698431365
transform -1 0 32704 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1022_
timestamp 1698431365
transform -1 0 31696 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1023_
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1024_
timestamp 1698431365
transform -1 0 31360 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1025_
timestamp 1698431365
transform -1 0 30464 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1026_
timestamp 1698431365
transform 1 0 29008 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1027_
timestamp 1698431365
transform -1 0 35168 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1028_
timestamp 1698431365
transform 1 0 30912 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1029_
timestamp 1698431365
transform 1 0 30800 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1030_
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1031_
timestamp 1698431365
transform 1 0 31808 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1032_
timestamp 1698431365
transform -1 0 34384 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1033_
timestamp 1698431365
transform -1 0 35840 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1034_
timestamp 1698431365
transform -1 0 34160 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1035_
timestamp 1698431365
transform -1 0 33264 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1036_
timestamp 1698431365
transform -1 0 34720 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1037_
timestamp 1698431365
transform 1 0 34608 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1038_
timestamp 1698431365
transform 1 0 31584 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1039_
timestamp 1698431365
transform 1 0 32032 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1040_
timestamp 1698431365
transform -1 0 33600 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1041_
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_4  _1042_
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1043_
timestamp 1698431365
transform 1 0 19936 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1044_
timestamp 1698431365
transform 1 0 23632 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1045_
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1046_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19488 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1047_
timestamp 1698431365
transform -1 0 25984 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1048_
timestamp 1698431365
transform -1 0 28784 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1049_
timestamp 1698431365
transform -1 0 34384 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1050_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37968 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1051_
timestamp 1698431365
transform 1 0 34832 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1052_
timestamp 1698431365
transform -1 0 34832 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1053_
timestamp 1698431365
transform 1 0 34048 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1054_
timestamp 1698431365
transform -1 0 35952 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1055_
timestamp 1698431365
transform 1 0 31808 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1056_
timestamp 1698431365
transform -1 0 31808 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1057_
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1058_
timestamp 1698431365
transform -1 0 28784 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1059_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25536 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1060_
timestamp 1698431365
transform -1 0 27888 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1061_
timestamp 1698431365
transform 1 0 26544 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1062_
timestamp 1698431365
transform 1 0 27664 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1063_
timestamp 1698431365
transform 1 0 32480 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1064_
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1065_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23744 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1066_
timestamp 1698431365
transform 1 0 33824 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1067_
timestamp 1698431365
transform 1 0 30240 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1068_
timestamp 1698431365
transform 1 0 30688 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1069_
timestamp 1698431365
transform -1 0 30688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1070_
timestamp 1698431365
transform 1 0 27552 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1071_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1072_
timestamp 1698431365
transform -1 0 26656 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1073_
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1074_
timestamp 1698431365
transform 1 0 29456 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1075_
timestamp 1698431365
transform -1 0 27552 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1076_
timestamp 1698431365
transform -1 0 26656 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1077_
timestamp 1698431365
transform 1 0 27664 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1078_
timestamp 1698431365
transform -1 0 27552 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1079_
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1080_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27104 0 1 10976
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1081_
timestamp 1698431365
transform -1 0 27328 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1082_
timestamp 1698431365
transform 1 0 24640 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1083_
timestamp 1698431365
transform 1 0 28112 0 -1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1084_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28336 0 -1 12544
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1085_
timestamp 1698431365
transform -1 0 30128 0 -1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1086_
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1087_
timestamp 1698431365
transform 1 0 30240 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1088_
timestamp 1698431365
transform 1 0 31808 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1089_
timestamp 1698431365
transform 1 0 34048 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1090_
timestamp 1698431365
transform -1 0 31808 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1091_
timestamp 1698431365
transform 1 0 34384 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1092_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31472 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1093_
timestamp 1698431365
transform -1 0 33824 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1094_
timestamp 1698431365
transform -1 0 34944 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1095_
timestamp 1698431365
transform -1 0 32704 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1096_
timestamp 1698431365
transform -1 0 34272 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1097_
timestamp 1698431365
transform -1 0 32704 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1098_
timestamp 1698431365
transform 1 0 33152 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1099_
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1100_
timestamp 1698431365
transform 1 0 32368 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1101_
timestamp 1698431365
transform -1 0 34048 0 1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1102_
timestamp 1698431365
transform -1 0 36400 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1103_
timestamp 1698431365
transform 1 0 34944 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1104_
timestamp 1698431365
transform -1 0 31696 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1105_
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1106_
timestamp 1698431365
transform 1 0 29904 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1107_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1108_
timestamp 1698431365
transform 1 0 28784 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1109_
timestamp 1698431365
transform -1 0 36512 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1110_
timestamp 1698431365
transform 1 0 33936 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1111_
timestamp 1698431365
transform 1 0 6944 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1112_
timestamp 1698431365
transform -1 0 20944 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1114_
timestamp 1698431365
transform 1 0 20160 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1115_
timestamp 1698431365
transform -1 0 20944 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1116_
timestamp 1698431365
transform -1 0 19600 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1117_
timestamp 1698431365
transform -1 0 20944 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1118_
timestamp 1698431365
transform -1 0 19600 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1119_
timestamp 1698431365
transform -1 0 18144 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1120_
timestamp 1698431365
transform 1 0 17360 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1121_
timestamp 1698431365
transform 1 0 21952 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _1122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21728 0 1 12544
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1123_
timestamp 1698431365
transform -1 0 32816 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1124_
timestamp 1698431365
transform 1 0 31808 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1125_
timestamp 1698431365
transform -1 0 33824 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1126_
timestamp 1698431365
transform 1 0 34384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1127_
timestamp 1698431365
transform 1 0 30352 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1128_
timestamp 1698431365
transform 1 0 31360 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1129_
timestamp 1698431365
transform 1 0 26656 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1130_
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1131_
timestamp 1698431365
transform -1 0 27664 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1132_
timestamp 1698431365
transform 1 0 27664 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1133_
timestamp 1698431365
transform 1 0 13776 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1134_
timestamp 1698431365
transform 1 0 14336 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23408 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1136_
timestamp 1698431365
transform 1 0 25312 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1137_
timestamp 1698431365
transform 1 0 26208 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1138_
timestamp 1698431365
transform 1 0 37520 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1139_
timestamp 1698431365
transform -1 0 38864 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1140_
timestamp 1698431365
transform -1 0 36064 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1141_
timestamp 1698431365
transform -1 0 32144 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1142_
timestamp 1698431365
transform -1 0 28224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1143_
timestamp 1698431365
transform -1 0 38528 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1144_
timestamp 1698431365
transform 1 0 37408 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1145_
timestamp 1698431365
transform -1 0 36960 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1146_
timestamp 1698431365
transform 1 0 29344 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1147_
timestamp 1698431365
transform 1 0 27104 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1148_
timestamp 1698431365
transform 1 0 22400 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1149_
timestamp 1698431365
transform -1 0 23856 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1150_
timestamp 1698431365
transform 1 0 19152 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1151_
timestamp 1698431365
transform 1 0 23632 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1152_
timestamp 1698431365
transform -1 0 18256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1153_
timestamp 1698431365
transform -1 0 21616 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1154_
timestamp 1698431365
transform -1 0 14672 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1155_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1156_
timestamp 1698431365
transform -1 0 5040 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1157_
timestamp 1698431365
transform -1 0 5264 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1158_
timestamp 1698431365
transform -1 0 5264 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1159_
timestamp 1698431365
transform -1 0 23520 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1160_
timestamp 1698431365
transform -1 0 15008 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1161_
timestamp 1698431365
transform -1 0 7840 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1162_
timestamp 1698431365
transform -1 0 6048 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1163_
timestamp 1698431365
transform -1 0 7280 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1164_
timestamp 1698431365
transform -1 0 13104 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1165_
timestamp 1698431365
transform -1 0 20720 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1166_
timestamp 1698431365
transform 1 0 13776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1167_
timestamp 1698431365
transform 1 0 15792 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1168_
timestamp 1698431365
transform 1 0 21616 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1169_
timestamp 1698431365
transform -1 0 23184 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1170_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1171_
timestamp 1698431365
transform -1 0 26880 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1172_
timestamp 1698431365
transform 1 0 28672 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1173_
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1174_
timestamp 1698431365
transform 1 0 34160 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1175_
timestamp 1698431365
transform 1 0 30688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1176_
timestamp 1698431365
transform -1 0 37296 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1177_
timestamp 1698431365
transform -1 0 31024 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1178_
timestamp 1698431365
transform -1 0 34832 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1179_
timestamp 1698431365
transform 1 0 35952 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1180_
timestamp 1698431365
transform 1 0 29232 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1181_
timestamp 1698431365
transform -1 0 26208 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1182_
timestamp 1698431365
transform 1 0 26656 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1183_
timestamp 1698431365
transform -1 0 24752 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1184_
timestamp 1698431365
transform -1 0 18256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1185_
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1186_
timestamp 1698431365
transform -1 0 12208 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1187_
timestamp 1698431365
transform 1 0 11088 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1188_
timestamp 1698431365
transform -1 0 14672 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1189_
timestamp 1698431365
transform -1 0 13328 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1190_
timestamp 1698431365
transform -1 0 21616 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1191_
timestamp 1698431365
transform -1 0 21616 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1192_
timestamp 1698431365
transform 1 0 19488 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1193_
timestamp 1698431365
transform -1 0 19040 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1194_
timestamp 1698431365
transform -1 0 11536 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1195_
timestamp 1698431365
transform 1 0 9184 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1196_
timestamp 1698431365
transform -1 0 7168 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1197_
timestamp 1698431365
transform -1 0 6832 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1198_
timestamp 1698431365
transform -1 0 5600 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1199_
timestamp 1698431365
transform 1 0 7280 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1200_
timestamp 1698431365
transform -1 0 8624 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1201_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13776 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1202_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13552 0 -1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1203_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34832 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1204_
timestamp 1698431365
transform 1 0 34608 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _1205_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32592 0 1 7840
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _1206_
timestamp 1698431365
transform -1 0 31696 0 -1 7840
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1207_
timestamp 1698431365
transform 1 0 23744 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1208_
timestamp 1698431365
transform 1 0 34272 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1209_
timestamp 1698431365
transform 1 0 34720 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1210_
timestamp 1698431365
transform 1 0 32816 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1211_
timestamp 1698431365
transform 1 0 27552 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1212_
timestamp 1698431365
transform 1 0 24528 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1213_
timestamp 1698431365
transform 1 0 20272 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1214_
timestamp 1698431365
transform 1 0 16576 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _1215_
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1216_
timestamp 1698431365
transform 1 0 14672 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1217_
timestamp 1698431365
transform 1 0 17136 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1218_
timestamp 1698431365
transform 1 0 10416 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1219_
timestamp 1698431365
transform 1 0 6608 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1220_
timestamp 1698431365
transform -1 0 5376 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1221_
timestamp 1698431365
transform 1 0 1904 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1222_
timestamp 1698431365
transform -1 0 6608 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _1223_
timestamp 1698431365
transform 1 0 11648 0 -1 28224
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1224_
timestamp 1698431365
transform 1 0 3584 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1225_
timestamp 1698431365
transform -1 0 6272 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1226_
timestamp 1698431365
transform 1 0 3696 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1227_
timestamp 1698431365
transform 1 0 8848 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1228_
timestamp 1698431365
transform 1 0 16464 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1229_
timestamp 1698431365
transform 1 0 11424 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1230_
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1231_
timestamp 1698431365
transform 1 0 18816 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1232_
timestamp 1698431365
transform 1 0 19488 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1233_
timestamp 1698431365
transform 1 0 23520 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1234_
timestamp 1698431365
transform 1 0 25872 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1235_
timestamp 1698431365
transform 1 0 22960 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1236_
timestamp 1698431365
transform 1 0 32816 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1237_
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1238_
timestamp 1698431365
transform 1 0 33712 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _1239_
timestamp 1698431365
transform 1 0 26544 0 -1 28224
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1240_
timestamp 1698431365
transform 1 0 29680 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1241_
timestamp 1698431365
transform 1 0 33488 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1242_
timestamp 1698431365
transform 1 0 26544 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1243_
timestamp 1698431365
transform 1 0 21952 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1244_
timestamp 1698431365
transform 1 0 23968 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _1245_
timestamp 1698431365
transform 1 0 21280 0 1 15680
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _1246_
timestamp 1698431365
transform 1 0 14784 0 1 14112
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1247_
timestamp 1698431365
transform 1 0 14448 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1248_
timestamp 1698431365
transform -1 0 13776 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _1249_
timestamp 1698431365
transform 1 0 18144 0 -1 9408
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_4  _1250_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18144 0 -1 7840
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_4  _1251_
timestamp 1698431365
transform 1 0 18032 0 -1 10976
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1252_
timestamp 1698431365
transform 1 0 14896 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1253_
timestamp 1698431365
transform 1 0 9856 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1254_
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1255_
timestamp 1698431365
transform 1 0 5040 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1256_
timestamp 1698431365
transform 1 0 2016 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1257_
timestamp 1698431365
transform -1 0 9184 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1258_
timestamp 1698431365
transform 1 0 7840 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0605__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0606__A2
timestamp 1698431365
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0607__A2
timestamp 1698431365
transform 1 0 16240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0609__A2
timestamp 1698431365
transform 1 0 17808 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0610__A2
timestamp 1698431365
transform 1 0 16352 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0612__A1
timestamp 1698431365
transform 1 0 19152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0612__A2
timestamp 1698431365
transform -1 0 21504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0613__A2
timestamp 1698431365
transform -1 0 21728 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0614__I
timestamp 1698431365
transform 1 0 27776 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0615__A2
timestamp 1698431365
transform -1 0 29792 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0616__A2
timestamp 1698431365
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0618__I0
timestamp 1698431365
transform -1 0 26992 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0618__S
timestamp 1698431365
transform -1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0621__I0
timestamp 1698431365
transform 1 0 31136 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0621__S
timestamp 1698431365
transform 1 0 31920 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0623__I
timestamp 1698431365
transform 1 0 35504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0624__A2
timestamp 1698431365
transform 1 0 35504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0625__A2
timestamp 1698431365
transform 1 0 35056 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0627__A2
timestamp 1698431365
transform 1 0 35504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0628__A2
timestamp 1698431365
transform 1 0 35056 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0670__A1
timestamp 1698431365
transform 1 0 4144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0677__I
timestamp 1698431365
transform -1 0 16352 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0678__I
timestamp 1698431365
transform -1 0 14672 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0680__A1
timestamp 1698431365
transform -1 0 18816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0680__B2
timestamp 1698431365
transform -1 0 19936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0687__I
timestamp 1698431365
transform 1 0 27440 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0689__I
timestamp 1698431365
transform -1 0 19376 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0694__A1
timestamp 1698431365
transform 1 0 28784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0696__A1
timestamp 1698431365
transform 1 0 31024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0696__C
timestamp 1698431365
transform 1 0 35840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0698__A1
timestamp 1698431365
transform 1 0 35952 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0700__A1
timestamp 1698431365
transform 1 0 35392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0701__A1
timestamp 1698431365
transform 1 0 31360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0704__A1
timestamp 1698431365
transform 1 0 29792 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0719__A1
timestamp 1698431365
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0726__A1
timestamp 1698431365
transform 1 0 5152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0729__A1
timestamp 1698431365
transform 1 0 7504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0780__A1
timestamp 1698431365
transform -1 0 31360 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0788__A1
timestamp 1698431365
transform 1 0 29232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0788__A3
timestamp 1698431365
transform -1 0 32592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0789__A1
timestamp 1698431365
transform 1 0 28000 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0790__A1
timestamp 1698431365
transform 1 0 26656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0790__A2
timestamp 1698431365
transform -1 0 24304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0791__A1
timestamp 1698431365
transform 1 0 12656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0792__A1
timestamp 1698431365
transform 1 0 9744 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0804__A1
timestamp 1698431365
transform 1 0 30688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0804__B1
timestamp 1698431365
transform -1 0 30464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0807__A1
timestamp 1698431365
transform 1 0 18368 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0807__A2
timestamp 1698431365
transform -1 0 19040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0809__I1
timestamp 1698431365
transform 1 0 33376 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0809__S
timestamp 1698431365
transform 1 0 27440 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0813__A1
timestamp 1698431365
transform 1 0 29792 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0815__A1
timestamp 1698431365
transform 1 0 35840 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0816__S
timestamp 1698431365
transform 1 0 34720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0819__I
timestamp 1698431365
transform 1 0 18928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0820__I
timestamp 1698431365
transform 1 0 22736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0825__I
timestamp 1698431365
transform 1 0 30352 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0826__A1
timestamp 1698431365
transform 1 0 29344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0826__B2
timestamp 1698431365
transform 1 0 29792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__I
timestamp 1698431365
transform 1 0 25872 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0828__A2
timestamp 1698431365
transform 1 0 33600 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0829__A1
timestamp 1698431365
transform 1 0 30240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0830__I
timestamp 1698431365
transform 1 0 26320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0833__A1
timestamp 1698431365
transform -1 0 31024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0833__B2
timestamp 1698431365
transform 1 0 33936 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0834__A2
timestamp 1698431365
transform 1 0 34832 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0835__A1
timestamp 1698431365
transform 1 0 33712 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0841__A1
timestamp 1698431365
transform 1 0 26992 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0841__B2
timestamp 1698431365
transform 1 0 26320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__S
timestamp 1698431365
transform -1 0 25088 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0846__A1
timestamp 1698431365
transform -1 0 29456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0846__B2
timestamp 1698431365
transform 1 0 26544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0847__A2
timestamp 1698431365
transform 1 0 29680 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0848__A1
timestamp 1698431365
transform 1 0 29344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0853__A1
timestamp 1698431365
transform 1 0 25200 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0853__B2
timestamp 1698431365
transform 1 0 25648 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0854__A2
timestamp 1698431365
transform -1 0 29792 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0855__A1
timestamp 1698431365
transform 1 0 26096 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0858__A1
timestamp 1698431365
transform 1 0 20272 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0858__B2
timestamp 1698431365
transform 1 0 24192 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0859__A2
timestamp 1698431365
transform 1 0 20720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0860__A1
timestamp 1698431365
transform 1 0 19824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0872__A1
timestamp 1698431365
transform 1 0 20944 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0872__B2
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0874__A2
timestamp 1698431365
transform 1 0 19936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__A1
timestamp 1698431365
transform 1 0 19040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0878__A1
timestamp 1698431365
transform 1 0 18368 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0878__B2
timestamp 1698431365
transform 1 0 17696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0879__S
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0886__A1
timestamp 1698431365
transform -1 0 20048 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0887__A1
timestamp 1698431365
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0888__S
timestamp 1698431365
transform -1 0 14896 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0892__A1
timestamp 1698431365
transform -1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0893__A1
timestamp 1698431365
transform 1 0 16352 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__A2
timestamp 1698431365
transform 1 0 19488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0895__A1
timestamp 1698431365
transform -1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0896__I
timestamp 1698431365
transform 1 0 22512 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0902__A1
timestamp 1698431365
transform -1 0 10640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0902__B2
timestamp 1698431365
transform 1 0 9968 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__A2
timestamp 1698431365
transform 1 0 12432 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0904__A1
timestamp 1698431365
transform -1 0 11088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0905__I
timestamp 1698431365
transform 1 0 19376 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0909__A1
timestamp 1698431365
transform 1 0 11424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0911__A1
timestamp 1698431365
transform -1 0 7952 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__A2
timestamp 1698431365
transform 1 0 7952 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0913__A1
timestamp 1698431365
transform 1 0 6832 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0918__A1
timestamp 1698431365
transform -1 0 6160 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0918__B2
timestamp 1698431365
transform -1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__A2
timestamp 1698431365
transform 1 0 6832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0920__A1
timestamp 1698431365
transform 1 0 5264 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__A1
timestamp 1698431365
transform 1 0 11424 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__B2
timestamp 1698431365
transform 1 0 11872 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__A2
timestamp 1698431365
transform 1 0 7056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0925__A1
timestamp 1698431365
transform 1 0 6608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0933__A1
timestamp 1698431365
transform -1 0 10304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__A1
timestamp 1698431365
transform 1 0 12432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0935__A2
timestamp 1698431365
transform 1 0 15792 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0936__A1
timestamp 1698431365
transform 1 0 11424 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0939__A1
timestamp 1698431365
transform 1 0 9632 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0939__B2
timestamp 1698431365
transform 1 0 8400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0940__A2
timestamp 1698431365
transform 1 0 6944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__A1
timestamp 1698431365
transform 1 0 6384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0943__B
timestamp 1698431365
transform -1 0 6048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0948__A1
timestamp 1698431365
transform 1 0 9296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0948__B2
timestamp 1698431365
transform 1 0 10864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0949__A2
timestamp 1698431365
transform -1 0 6272 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0950__A1
timestamp 1698431365
transform 1 0 4704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0953__A1
timestamp 1698431365
transform 1 0 10416 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0954__A1
timestamp 1698431365
transform 1 0 10976 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0955__A2
timestamp 1698431365
transform 1 0 6720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0956__A1
timestamp 1698431365
transform -1 0 4368 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0963__A1
timestamp 1698431365
transform 1 0 10192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0963__B2
timestamp 1698431365
transform 1 0 7952 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0964__A2
timestamp 1698431365
transform -1 0 10192 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0965__A1
timestamp 1698431365
transform 1 0 8512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0966__A1
timestamp 1698431365
transform 1 0 12208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__A1
timestamp 1698431365
transform 1 0 14896 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0969__A1
timestamp 1698431365
transform 1 0 15344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0971__A2
timestamp 1698431365
transform -1 0 14896 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0972__A1
timestamp 1698431365
transform -1 0 12320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0973__A1
timestamp 1698431365
transform 1 0 19712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0975__A1
timestamp 1698431365
transform 1 0 19264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0979__A1
timestamp 1698431365
transform -1 0 17808 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0979__B2
timestamp 1698431365
transform -1 0 18144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__A1
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__A2
timestamp 1698431365
transform 1 0 17472 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0981__A1
timestamp 1698431365
transform 1 0 17024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0982__A1
timestamp 1698431365
transform -1 0 14224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0983__A1
timestamp 1698431365
transform 1 0 19264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__B2
timestamp 1698431365
transform -1 0 18368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__A1
timestamp 1698431365
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__A2
timestamp 1698431365
transform 1 0 16352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0987__A1
timestamp 1698431365
transform 1 0 18368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0989__A1
timestamp 1698431365
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__A1
timestamp 1698431365
transform 1 0 24192 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__B2
timestamp 1698431365
transform 1 0 23744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0996__A2
timestamp 1698431365
transform 1 0 24304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0997__A1
timestamp 1698431365
transform 1 0 25312 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__A1
timestamp 1698431365
transform 1 0 20160 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0999__A1
timestamp 1698431365
transform 1 0 20272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1001__A1
timestamp 1698431365
transform 1 0 19600 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A2
timestamp 1698431365
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1004__A1
timestamp 1698431365
transform 1 0 19376 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1007__A1
timestamp 1698431365
transform 1 0 28448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1008__A1
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__A1
timestamp 1698431365
transform 1 0 27328 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1010__S
timestamp 1698431365
transform -1 0 23856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1013__A1
timestamp 1698431365
transform 1 0 27888 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1014__A1
timestamp 1698431365
transform 1 0 28112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1015__B2
timestamp 1698431365
transform -1 0 27216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__A2
timestamp 1698431365
transform 1 0 25424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__A1
timestamp 1698431365
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1020__A1
timestamp 1698431365
transform -1 0 33152 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1022__A1
timestamp 1698431365
transform 1 0 31920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1022__A2
timestamp 1698431365
transform 1 0 31696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__A1
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1024__A1
timestamp 1698431365
transform 1 0 30240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__A1
timestamp 1698431365
transform 1 0 31136 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__C
timestamp 1698431365
transform 1 0 31584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1026__A2
timestamp 1698431365
transform 1 0 30912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1028__A1
timestamp 1698431365
transform 1 0 32144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1028__B
timestamp 1698431365
transform 1 0 30688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1030__A1
timestamp 1698431365
transform 1 0 34272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1030__B2
timestamp 1698431365
transform 1 0 34832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1030__C
timestamp 1698431365
transform 1 0 35280 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1031__A2
timestamp 1698431365
transform 1 0 34384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1034__A1
timestamp 1698431365
transform 1 0 35392 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__A1
timestamp 1698431365
transform 1 0 32032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1036__S
timestamp 1698431365
transform 1 0 35504 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__A2
timestamp 1698431365
transform 1 0 31920 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A2
timestamp 1698431365
transform 1 0 32256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__B
timestamp 1698431365
transform 1 0 34944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1041__A2
timestamp 1698431365
transform 1 0 35840 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__A1
timestamp 1698431365
transform 1 0 31360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__A1
timestamp 1698431365
transform 1 0 35056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1051__A1
timestamp 1698431365
transform 1 0 35952 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__A1
timestamp 1698431365
transform 1 0 35504 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__A1
timestamp 1698431365
transform -1 0 32256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__A1
timestamp 1698431365
transform 1 0 30576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1059__A1
timestamp 1698431365
transform 1 0 30128 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__A1
timestamp 1698431365
transform -1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A1
timestamp 1698431365
transform 1 0 31584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__A1
timestamp 1698431365
transform 1 0 29232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__A1
timestamp 1698431365
transform 1 0 30912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__A1
timestamp 1698431365
transform 1 0 30912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1088__A1
timestamp 1698431365
transform -1 0 31808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__A1
timestamp 1698431365
transform -1 0 31248 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__A1
timestamp 1698431365
transform 1 0 35616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__A1
timestamp 1698431365
transform -1 0 35392 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1104__A1
timestamp 1698431365
transform 1 0 31920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__I
timestamp 1698431365
transform -1 0 28000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1138__I
timestamp 1698431365
transform 1 0 37296 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__I
timestamp 1698431365
transform 1 0 39088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1140__I
timestamp 1698431365
transform 1 0 35392 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1141__I
timestamp 1698431365
transform 1 0 32368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1142__I
timestamp 1698431365
transform 1 0 27440 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1143__I
timestamp 1698431365
transform 1 0 37856 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1144__I
timestamp 1698431365
transform 1 0 37184 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1145__I
timestamp 1698431365
transform 1 0 37184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1146__I
timestamp 1698431365
transform 1 0 30576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1147__I
timestamp 1698431365
transform -1 0 28560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__I
timestamp 1698431365
transform 1 0 24080 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1150__I
timestamp 1698431365
transform -1 0 20048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1151__I
timestamp 1698431365
transform 1 0 24304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__I
timestamp 1698431365
transform 1 0 18704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__I
timestamp 1698431365
transform 1 0 22400 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1154__I
timestamp 1698431365
transform -1 0 14784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__I
timestamp 1698431365
transform 1 0 10080 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1156__I
timestamp 1698431365
transform 1 0 5712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1157__I
timestamp 1698431365
transform -1 0 4816 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__I
timestamp 1698431365
transform -1 0 4816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1160__I
timestamp 1698431365
transform 1 0 15232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1161__I
timestamp 1698431365
transform 1 0 8064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__I
timestamp 1698431365
transform 1 0 6048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1163__I
timestamp 1698431365
transform 1 0 7280 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1164__I
timestamp 1698431365
transform 1 0 11200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__I
timestamp 1698431365
transform 1 0 18592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1166__I
timestamp 1698431365
transform 1 0 13552 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1167__I
timestamp 1698431365
transform 1 0 16464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1168__I
timestamp 1698431365
transform 1 0 21392 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1169__I
timestamp 1698431365
transform 1 0 23968 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1171__I
timestamp 1698431365
transform 1 0 27888 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1172__I
timestamp 1698431365
transform 1 0 30240 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1173__I
timestamp 1698431365
transform 1 0 25760 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1174__I
timestamp 1698431365
transform 1 0 34384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1175__I
timestamp 1698431365
transform -1 0 33376 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1176__I
timestamp 1698431365
transform 1 0 37520 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1177__I
timestamp 1698431365
transform 1 0 32032 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1178__I
timestamp 1698431365
transform 1 0 35952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1179__I
timestamp 1698431365
transform -1 0 36176 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1180__I
timestamp 1698431365
transform 1 0 30016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1181__I
timestamp 1698431365
transform 1 0 26208 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1182__I
timestamp 1698431365
transform 1 0 28224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1183__I
timestamp 1698431365
transform 1 0 28000 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1184__I
timestamp 1698431365
transform 1 0 19040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1185__I
timestamp 1698431365
transform -1 0 15456 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1190__I
timestamp 1698431365
transform -1 0 22064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1191__I
timestamp 1698431365
transform -1 0 22512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__I
timestamp 1698431365
transform 1 0 19264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__I
timestamp 1698431365
transform 1 0 19264 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1201__CLK
timestamp 1698431365
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1202__CLK
timestamp 1698431365
transform -1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1203__CLK
timestamp 1698431365
transform 1 0 36064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1204__CLK
timestamp 1698431365
transform 1 0 34608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1205__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1206__CLK
timestamp 1698431365
transform -1 0 31920 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1207__CLK
timestamp 1698431365
transform -1 0 28448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1208__CLK
timestamp 1698431365
transform 1 0 36064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1209__CLK
timestamp 1698431365
transform 1 0 35056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__CLK
timestamp 1698431365
transform 1 0 33824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1211__CLK
timestamp 1698431365
transform -1 0 31696 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1212__CLK
timestamp 1698431365
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1213__CLK
timestamp 1698431365
transform 1 0 27552 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1214__CLK
timestamp 1698431365
transform 1 0 16352 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1215__CLK
timestamp 1698431365
transform 1 0 25424 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__CLK
timestamp 1698431365
transform 1 0 14448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1217__CLK
timestamp 1698431365
transform 1 0 16576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1218__CLK
timestamp 1698431365
transform 1 0 14112 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1219__CLK
timestamp 1698431365
transform 1 0 10640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1220__CLK
timestamp 1698431365
transform 1 0 5376 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1221__CLK
timestamp 1698431365
transform 1 0 6496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1222__CLK
timestamp 1698431365
transform 1 0 6832 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1223__CLK
timestamp 1698431365
transform 1 0 15904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1224__CLK
timestamp 1698431365
transform 1 0 7392 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1225__CLK
timestamp 1698431365
transform 1 0 6272 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1226__CLK
timestamp 1698431365
transform 1 0 7504 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1227__CLK
timestamp 1698431365
transform 1 0 10752 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1228__CLK
timestamp 1698431365
transform -1 0 15344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1229__CLK
timestamp 1698431365
transform 1 0 13104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1230__CLK
timestamp 1698431365
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1231__CLK
timestamp 1698431365
transform 1 0 22624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1232__CLK
timestamp 1698431365
transform -1 0 19264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1233__CLK
timestamp 1698431365
transform 1 0 29792 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1234__CLK
timestamp 1698431365
transform -1 0 31360 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1235__CLK
timestamp 1698431365
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1236__CLK
timestamp 1698431365
transform 1 0 34048 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1237__CLK
timestamp 1698431365
transform 1 0 34496 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1238__CLK
timestamp 1698431365
transform 1 0 35168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1239__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1240__CLK
timestamp 1698431365
transform 1 0 35504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1241__CLK
timestamp 1698431365
transform 1 0 35056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1242__CLK
timestamp 1698431365
transform 1 0 31472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1243__CLK
timestamp 1698431365
transform 1 0 25760 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1244__CLK
timestamp 1698431365
transform 1 0 29120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1245__CLK
timestamp 1698431365
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1246__CLK
timestamp 1698431365
transform 1 0 13664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1247__CLK
timestamp 1698431365
transform 1 0 14224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1248__CLK
timestamp 1698431365
transform 1 0 13664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1252__CLK
timestamp 1698431365
transform -1 0 15456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1253__CLK
timestamp 1698431365
transform -1 0 13776 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1254__CLK
timestamp 1698431365
transform -1 0 12656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__CLK
timestamp 1698431365
transform 1 0 8512 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1256__CLK
timestamp 1698431365
transform 1 0 4816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1257__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1258__CLK
timestamp 1698431365
transform 1 0 12432 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clock_I
timestamp 1698431365
transform -1 0 18704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_clock_I
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_clock_I
timestamp 1698431365
transform 1 0 15680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_clock_I
timestamp 1698431365
transform 1 0 28672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_clock_I
timestamp 1698431365
transform -1 0 25536 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 40432 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 1792 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 4032 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 2016 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 4032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 2464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 2688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 2464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 2464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 11088 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 39536 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 11536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 19376 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 18816 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 26208 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 28336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 31584 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 34944 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 39984 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform -1 0 39760 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 40208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 39760 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 39760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 26320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 39088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 20496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 38640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 3696 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 3584 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 23184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output64_I
timestamp 1698431365
transform 1 0 38640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output70_I
timestamp 1698431365
transform 1 0 3360 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output71_I
timestamp 1698431365
transform -1 0 3808 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clock dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18368 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clock
timestamp 1698431365
transform -1 0 16128 0 -1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clock
timestamp 1698431365
transform -1 0 15680 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clock
timestamp 1698431365
transform 1 0 27104 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clock
timestamp 1698431365
transform 1 0 26208 0 -1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_146 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_150 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18144 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_161
timestamp 1698431365
transform 1 0 19376 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698431365
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_180
timestamp 1698431365
transform 1 0 21504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_191 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_214
timestamp 1698431365
transform 1 0 25312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_233
timestamp 1698431365
transform 1 0 27440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698431365
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698431365
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_152
timestamp 1698431365
transform 1 0 18368 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_184 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21952 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_200
timestamp 1698431365
transform 1 0 23744 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_208
timestamp 1698431365
transform 1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_222
timestamp 1698431365
transform 1 0 26208 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_225
timestamp 1698431365
transform 1 0 26544 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_257
timestamp 1698431365
transform 1 0 30128 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_273
timestamp 1698431365
transform 1 0 31920 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_277
timestamp 1698431365
transform 1 0 32368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698431365
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698431365
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_181
timestamp 1698431365
transform 1 0 21616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_185
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_189
timestamp 1698431365
transform 1 0 22512 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_197
timestamp 1698431365
transform 1 0 23408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_199
timestamp 1698431365
transform 1 0 23632 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_234
timestamp 1698431365
transform 1 0 27552 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_238
timestamp 1698431365
transform 1 0 28000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_242
timestamp 1698431365
transform 1 0 28448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_244
timestamp 1698431365
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_263
timestamp 1698431365
transform 1 0 30800 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_273
timestamp 1698431365
transform 1 0 31920 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_305
timestamp 1698431365
transform 1 0 35504 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_313
timestamp 1698431365
transform 1 0 36400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_190
timestamp 1698431365
transform 1 0 22624 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_194
timestamp 1698431365
transform 1 0 23072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_202
timestamp 1698431365
transform 1 0 23968 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_220
timestamp 1698431365
transform 1 0 25984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_224
timestamp 1698431365
transform 1 0 26432 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_226
timestamp 1698431365
transform 1 0 26656 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_229
timestamp 1698431365
transform 1 0 26992 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_275
timestamp 1698431365
transform 1 0 32144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_286
timestamp 1698431365
transform 1 0 33376 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_302
timestamp 1698431365
transform 1 0 35168 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_310
timestamp 1698431365
transform 1 0 36064 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_342
timestamp 1698431365
transform 1 0 39648 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698431365
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_139
timestamp 1698431365
transform 1 0 16912 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_155
timestamp 1698431365
transform 1 0 18704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_181
timestamp 1698431365
transform 1 0 21616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_183
timestamp 1698431365
transform 1 0 21840 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_259
timestamp 1698431365
transform 1 0 30352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_263
timestamp 1698431365
transform 1 0 30800 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_267
timestamp 1698431365
transform 1 0 31248 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_269
timestamp 1698431365
transform 1 0 31472 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_272
timestamp 1698431365
transform 1 0 31808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_276
timestamp 1698431365
transform 1 0 32256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_278
timestamp 1698431365
transform 1 0 32480 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_200
timestamp 1698431365
transform 1 0 23744 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_237
timestamp 1698431365
transform 1 0 27888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_262
timestamp 1698431365
transform 1 0 30688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_266
timestamp 1698431365
transform 1 0 31136 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_295
timestamp 1698431365
transform 1 0 34384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_299
timestamp 1698431365
transform 1 0 34832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_303
timestamp 1698431365
transform 1 0 35280 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_335
timestamp 1698431365
transform 1 0 38864 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_343
timestamp 1698431365
transform 1 0 39760 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_347
timestamp 1698431365
transform 1 0 40208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_69
timestamp 1698431365
transform 1 0 9072 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_77
timestamp 1698431365
transform 1 0 9968 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_81
timestamp 1698431365
transform 1 0 10416 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_91
timestamp 1698431365
transform 1 0 11536 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_115
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_122
timestamp 1698431365
transform 1 0 15008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_126
timestamp 1698431365
transform 1 0 15456 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_158
timestamp 1698431365
transform 1 0 19040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_183
timestamp 1698431365
transform 1 0 21840 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_207
timestamp 1698431365
transform 1 0 24528 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_239
timestamp 1698431365
transform 1 0 28112 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_266
timestamp 1698431365
transform 1 0 31136 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_270
timestamp 1698431365
transform 1 0 31584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_300
timestamp 1698431365
transform 1 0 34944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_304
timestamp 1698431365
transform 1 0 35392 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_312
timestamp 1698431365
transform 1 0 36288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_107
timestamp 1698431365
transform 1 0 13328 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_189
timestamp 1698431365
transform 1 0 22512 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_205
timestamp 1698431365
transform 1 0 24304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_221
timestamp 1698431365
transform 1 0 26096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_223
timestamp 1698431365
transform 1 0 26320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_257
timestamp 1698431365
transform 1 0 30128 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_262
timestamp 1698431365
transform 1 0 30688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_266
timestamp 1698431365
transform 1 0 31136 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_294
timestamp 1698431365
transform 1 0 34272 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_296
timestamp 1698431365
transform 1 0 34496 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_335
timestamp 1698431365
transform 1 0 38864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_339
timestamp 1698431365
transform 1 0 39312 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_347
timestamp 1698431365
transform 1 0 40208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_45
timestamp 1698431365
transform 1 0 6384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_47
timestamp 1698431365
transform 1 0 6608 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_52
timestamp 1698431365
transform 1 0 7168 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_68
timestamp 1698431365
transform 1 0 8960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_119
timestamp 1698431365
transform 1 0 14672 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_155
timestamp 1698431365
transform 1 0 18704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_179
timestamp 1698431365
transform 1 0 21392 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_196
timestamp 1698431365
transform 1 0 23296 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_313
timestamp 1698431365
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_327
timestamp 1698431365
transform 1 0 37968 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_343
timestamp 1698431365
transform 1 0 39760 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_347
timestamp 1698431365
transform 1 0 40208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_18
timestamp 1698431365
transform 1 0 3360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_26
timestamp 1698431365
transform 1 0 4256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_30
timestamp 1698431365
transform 1 0 4704 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_62
timestamp 1698431365
transform 1 0 8288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_80
timestamp 1698431365
transform 1 0 10304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_158
timestamp 1698431365
transform 1 0 19040 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_238
timestamp 1698431365
transform 1 0 28000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_240
timestamp 1698431365
transform 1 0 28224 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_271
timestamp 1698431365
transform 1 0 31696 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_275
timestamp 1698431365
transform 1 0 32144 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_278
timestamp 1698431365
transform 1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_303
timestamp 1698431365
transform 1 0 35280 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_307
timestamp 1698431365
transform 1 0 35728 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_311
timestamp 1698431365
transform 1 0 36176 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_343
timestamp 1698431365
transform 1 0 39760 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_347
timestamp 1698431365
transform 1 0 40208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_49
timestamp 1698431365
transform 1 0 6832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_97
timestamp 1698431365
transform 1 0 12208 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_109
timestamp 1698431365
transform 1 0 13552 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_128
timestamp 1698431365
transform 1 0 15680 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_144
timestamp 1698431365
transform 1 0 17472 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_148
timestamp 1698431365
transform 1 0 17920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_179
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_260
timestamp 1698431365
transform 1 0 30464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_267
timestamp 1698431365
transform 1 0 31248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_271
timestamp 1698431365
transform 1 0 31696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_275
timestamp 1698431365
transform 1 0 32144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_289
timestamp 1698431365
transform 1 0 33712 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_327
timestamp 1698431365
transform 1 0 37968 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_331
timestamp 1698431365
transform 1 0 38416 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_335
timestamp 1698431365
transform 1 0 38864 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_18
timestamp 1698431365
transform 1 0 3360 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_26
timestamp 1698431365
transform 1 0 4256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_30
timestamp 1698431365
transform 1 0 4704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_38
timestamp 1698431365
transform 1 0 5600 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_40
timestamp 1698431365
transform 1 0 5824 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_76
timestamp 1698431365
transform 1 0 9856 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_80
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_132
timestamp 1698431365
transform 1 0 16128 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_146
timestamp 1698431365
transform 1 0 17696 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_149
timestamp 1698431365
transform 1 0 18032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_153
timestamp 1698431365
transform 1 0 18480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_155
timestamp 1698431365
transform 1 0 18704 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_165
timestamp 1698431365
transform 1 0 19824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_167
timestamp 1698431365
transform 1 0 20048 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_243
timestamp 1698431365
transform 1 0 28560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_268
timestamp 1698431365
transform 1 0 31360 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_333
timestamp 1698431365
transform 1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_65
timestamp 1698431365
transform 1 0 8624 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_97
timestamp 1698431365
transform 1 0 12208 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_109
timestamp 1698431365
transform 1 0 13552 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_112
timestamp 1698431365
transform 1 0 13888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_116
timestamp 1698431365
transform 1 0 14336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_156
timestamp 1698431365
transform 1 0 18816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_160
timestamp 1698431365
transform 1 0 19264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698431365
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_271
timestamp 1698431365
transform 1 0 31696 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_275
timestamp 1698431365
transform 1 0 32144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_277
timestamp 1698431365
transform 1 0 32368 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_288
timestamp 1698431365
transform 1 0 33600 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_304
timestamp 1698431365
transform 1 0 35392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_308
timestamp 1698431365
transform 1 0 35840 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_312
timestamp 1698431365
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_333
timestamp 1698431365
transform 1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_76
timestamp 1698431365
transform 1 0 9856 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_80
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_119
timestamp 1698431365
transform 1 0 14672 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_123
timestamp 1698431365
transform 1 0 15120 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_134
timestamp 1698431365
transform 1 0 16352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_151
timestamp 1698431365
transform 1 0 18256 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_198
timestamp 1698431365
transform 1 0 23520 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_224
timestamp 1698431365
transform 1 0 26432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_276
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_299
timestamp 1698431365
transform 1 0 34832 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_303
timestamp 1698431365
transform 1 0 35280 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_307
timestamp 1698431365
transform 1 0 35728 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_311
timestamp 1698431365
transform 1 0 36176 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_327
timestamp 1698431365
transform 1 0 37968 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_345
timestamp 1698431365
transform 1 0 39984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_16
timestamp 1698431365
transform 1 0 3136 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698431365
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_45
timestamp 1698431365
transform 1 0 6384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_81
timestamp 1698431365
transform 1 0 10416 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_85
timestamp 1698431365
transform 1 0 10864 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_93
timestamp 1698431365
transform 1 0 11760 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_95
timestamp 1698431365
transform 1 0 11984 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_111
timestamp 1698431365
transform 1 0 13776 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_151
timestamp 1698431365
transform 1 0 18256 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_233
timestamp 1698431365
transform 1 0 27440 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_241
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_262
timestamp 1698431365
transform 1 0 30688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_299
timestamp 1698431365
transform 1 0 34832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_303
timestamp 1698431365
transform 1 0 35280 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_307
timestamp 1698431365
transform 1 0 35728 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_313
timestamp 1698431365
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_333
timestamp 1698431365
transform 1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_16
timestamp 1698431365
transform 1 0 3136 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_48
timestamp 1698431365
transform 1 0 6720 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_64
timestamp 1698431365
transform 1 0 8512 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698431365
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_76
timestamp 1698431365
transform 1 0 9856 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_91
timestamp 1698431365
transform 1 0 11536 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_117
timestamp 1698431365
transform 1 0 14448 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_121
timestamp 1698431365
transform 1 0 14896 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_131
timestamp 1698431365
transform 1 0 16016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_135
timestamp 1698431365
transform 1 0 16464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_137
timestamp 1698431365
transform 1 0 16688 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_147
timestamp 1698431365
transform 1 0 17808 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_197
timestamp 1698431365
transform 1 0 23408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_201
timestamp 1698431365
transform 1 0 23856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_321
timestamp 1698431365
transform 1 0 37296 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_329
timestamp 1698431365
transform 1 0 38192 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_333
timestamp 1698431365
transform 1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_345
timestamp 1698431365
transform 1 0 39984 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_18
timestamp 1698431365
transform 1 0 3360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_22
timestamp 1698431365
transform 1 0 3808 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_26
timestamp 1698431365
transform 1 0 4256 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_28
timestamp 1698431365
transform 1 0 4480 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_41
timestamp 1698431365
transform 1 0 5936 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_44
timestamp 1698431365
transform 1 0 6272 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_48
timestamp 1698431365
transform 1 0 6720 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_74
timestamp 1698431365
transform 1 0 9632 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_102
timestamp 1698431365
transform 1 0 12768 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698431365
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_119
timestamp 1698431365
transform 1 0 14672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_123
timestamp 1698431365
transform 1 0 15120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_127
timestamp 1698431365
transform 1 0 15568 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_131
timestamp 1698431365
transform 1 0 16016 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_134
timestamp 1698431365
transform 1 0 16352 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_138
timestamp 1698431365
transform 1 0 16800 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_142
timestamp 1698431365
transform 1 0 17248 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_146
timestamp 1698431365
transform 1 0 17696 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_150
timestamp 1698431365
transform 1 0 18144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_154
timestamp 1698431365
transform 1 0 18592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698431365
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_187
timestamp 1698431365
transform 1 0 22288 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_236
timestamp 1698431365
transform 1 0 27776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_240
timestamp 1698431365
transform 1 0 28224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698431365
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_299
timestamp 1698431365
transform 1 0 34832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_303
timestamp 1698431365
transform 1 0 35280 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_307
timestamp 1698431365
transform 1 0 35728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_333
timestamp 1698431365
transform 1 0 38640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_4
timestamp 1698431365
transform 1 0 1792 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_39
timestamp 1698431365
transform 1 0 5712 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_41
timestamp 1698431365
transform 1 0 5936 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_46
timestamp 1698431365
transform 1 0 6496 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_53
timestamp 1698431365
transform 1 0 7280 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_57
timestamp 1698431365
transform 1 0 7728 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_84
timestamp 1698431365
transform 1 0 10752 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_117
timestamp 1698431365
transform 1 0 14448 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_119
timestamp 1698431365
transform 1 0 14672 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_136
timestamp 1698431365
transform 1 0 16576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_152
timestamp 1698431365
transform 1 0 18368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_156
timestamp 1698431365
transform 1 0 18816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_158
timestamp 1698431365
transform 1 0 19040 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_175
timestamp 1698431365
transform 1 0 20944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_177
timestamp 1698431365
transform 1 0 21168 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_186
timestamp 1698431365
transform 1 0 22176 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_190
timestamp 1698431365
transform 1 0 22624 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_201
timestamp 1698431365
transform 1 0 23856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_205
timestamp 1698431365
transform 1 0 24304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_230
timestamp 1698431365
transform 1 0 27104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_234
timestamp 1698431365
transform 1 0 27552 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_238
timestamp 1698431365
transform 1 0 28000 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_242
timestamp 1698431365
transform 1 0 28448 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_246
timestamp 1698431365
transform 1 0 28896 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_250
timestamp 1698431365
transform 1 0 29344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_254
timestamp 1698431365
transform 1 0 29792 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_258
timestamp 1698431365
transform 1 0 30240 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_264
timestamp 1698431365
transform 1 0 30912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_268
timestamp 1698431365
transform 1 0 31360 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_270
timestamp 1698431365
transform 1 0 31584 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_273
timestamp 1698431365
transform 1 0 31920 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698431365
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_299
timestamp 1698431365
transform 1 0 34832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_303
timestamp 1698431365
transform 1 0 35280 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_307
timestamp 1698431365
transform 1 0 35728 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_339
timestamp 1698431365
transform 1 0 39312 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_347
timestamp 1698431365
transform 1 0 40208 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_22
timestamp 1698431365
transform 1 0 3808 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_24
timestamp 1698431365
transform 1 0 4032 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_60
timestamp 1698431365
transform 1 0 8064 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_69
timestamp 1698431365
transform 1 0 9072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698431365
transform 1 0 9520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_77
timestamp 1698431365
transform 1 0 9968 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_81
timestamp 1698431365
transform 1 0 10416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_132
timestamp 1698431365
transform 1 0 16128 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_181
timestamp 1698431365
transform 1 0 21616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_183
timestamp 1698431365
transform 1 0 21840 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_219
timestamp 1698431365
transform 1 0 25872 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_228
timestamp 1698431365
transform 1 0 26880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_230
timestamp 1698431365
transform 1 0 27104 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_251
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_253
timestamp 1698431365
transform 1 0 29680 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_272
timestamp 1698431365
transform 1 0 31808 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_276
timestamp 1698431365
transform 1 0 32256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_303
timestamp 1698431365
transform 1 0 35280 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_307
timestamp 1698431365
transform 1 0 35728 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698431365
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_319
timestamp 1698431365
transform 1 0 37072 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_326
timestamp 1698431365
transform 1 0 37856 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_334
timestamp 1698431365
transform 1 0 38752 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_338
timestamp 1698431365
transform 1 0 39200 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_340
timestamp 1698431365
transform 1 0 39424 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_16
timestamp 1698431365
transform 1 0 3136 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_22
timestamp 1698431365
transform 1 0 3808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_26
timestamp 1698431365
transform 1 0 4256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_32
timestamp 1698431365
transform 1 0 4928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_83
timestamp 1698431365
transform 1 0 10640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_87
timestamp 1698431365
transform 1 0 11088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_95
timestamp 1698431365
transform 1 0 11984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_99
timestamp 1698431365
transform 1 0 12432 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_151
timestamp 1698431365
transform 1 0 18256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_232
timestamp 1698431365
transform 1 0 27328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_236
timestamp 1698431365
transform 1 0 27776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_240
timestamp 1698431365
transform 1 0 28224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_244
timestamp 1698431365
transform 1 0 28672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_246
timestamp 1698431365
transform 1 0 28896 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_271
timestamp 1698431365
transform 1 0 31696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_275
timestamp 1698431365
transform 1 0 32144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_332
timestamp 1698431365
transform 1 0 38528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_334
timestamp 1698431365
transform 1 0 38752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_18
timestamp 1698431365
transform 1 0 3360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_20
timestamp 1698431365
transform 1 0 3584 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_23
timestamp 1698431365
transform 1 0 3920 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_39
timestamp 1698431365
transform 1 0 5712 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_70
timestamp 1698431365
transform 1 0 9184 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_72
timestamp 1698431365
transform 1 0 9408 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_86
timestamp 1698431365
transform 1 0 10976 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_90
timestamp 1698431365
transform 1 0 11424 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_103
timestamp 1698431365
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_158
timestamp 1698431365
transform 1 0 19040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_162
timestamp 1698431365
transform 1 0 19488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_166
timestamp 1698431365
transform 1 0 19936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_224
timestamp 1698431365
transform 1 0 26432 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_237
timestamp 1698431365
transform 1 0 27888 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_252
timestamp 1698431365
transform 1 0 29568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_256
timestamp 1698431365
transform 1 0 30016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_260
timestamp 1698431365
transform 1 0 30464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_262
timestamp 1698431365
transform 1 0 30688 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_271
timestamp 1698431365
transform 1 0 31696 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_308
timestamp 1698431365
transform 1 0 35840 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698431365
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_325
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_328
timestamp 1698431365
transform 1 0 38080 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_336
timestamp 1698431365
transform 1 0 38976 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_340
timestamp 1698431365
transform 1 0 39424 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_84
timestamp 1698431365
transform 1 0 10752 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_88
timestamp 1698431365
transform 1 0 11200 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_96
timestamp 1698431365
transform 1 0 12096 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_113
timestamp 1698431365
transform 1 0 14000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_148
timestamp 1698431365
transform 1 0 17920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698431365
transform 1 0 24528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_268
timestamp 1698431365
transform 1 0 31360 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_332
timestamp 1698431365
transform 1 0 38528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_334
timestamp 1698431365
transform 1 0 38752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_24
timestamp 1698431365
transform 1 0 4032 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_28
timestamp 1698431365
transform 1 0 4480 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_33
timestamp 1698431365
transform 1 0 5040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_41
timestamp 1698431365
transform 1 0 5936 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_46
timestamp 1698431365
transform 1 0 6496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_50
timestamp 1698431365
transform 1 0 6944 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_57
timestamp 1698431365
transform 1 0 7728 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_79
timestamp 1698431365
transform 1 0 10192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_83
timestamp 1698431365
transform 1 0 10640 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_111
timestamp 1698431365
transform 1 0 13776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_115
timestamp 1698431365
transform 1 0 14224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_119
timestamp 1698431365
transform 1 0 14672 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_123
timestamp 1698431365
transform 1 0 15120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_125
timestamp 1698431365
transform 1 0 15344 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_147
timestamp 1698431365
transform 1 0 17808 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_158
timestamp 1698431365
transform 1 0 19040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_162
timestamp 1698431365
transform 1 0 19488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_166
timestamp 1698431365
transform 1 0 19936 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_168
timestamp 1698431365
transform 1 0 20160 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_190
timestamp 1698431365
transform 1 0 22624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_227
timestamp 1698431365
transform 1 0 26768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_231
timestamp 1698431365
transform 1 0 27216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_235
timestamp 1698431365
transform 1 0 27664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_239
timestamp 1698431365
transform 1 0 28112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_259
timestamp 1698431365
transform 1 0 30352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_263
timestamp 1698431365
transform 1 0 30800 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_267
timestamp 1698431365
transform 1 0 31248 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_271
timestamp 1698431365
transform 1 0 31696 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_275
timestamp 1698431365
transform 1 0 32144 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_278
timestamp 1698431365
transform 1 0 32480 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_298
timestamp 1698431365
transform 1 0 34720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_302
timestamp 1698431365
transform 1 0 35168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_306
timestamp 1698431365
transform 1 0 35616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_310
timestamp 1698431365
transform 1 0 36064 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_333
timestamp 1698431365
transform 1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_16
timestamp 1698431365
transform 1 0 3136 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_20
timestamp 1698431365
transform 1 0 3584 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_38
timestamp 1698431365
transform 1 0 5600 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_46
timestamp 1698431365
transform 1 0 6496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_50
timestamp 1698431365
transform 1 0 6944 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_109
timestamp 1698431365
transform 1 0 13552 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_125
timestamp 1698431365
transform 1 0 15344 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_129
timestamp 1698431365
transform 1 0 15792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_150
timestamp 1698431365
transform 1 0 18144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_154
timestamp 1698431365
transform 1 0 18592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_158
timestamp 1698431365
transform 1 0 19040 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_161
timestamp 1698431365
transform 1 0 19376 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_195
timestamp 1698431365
transform 1 0 23184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_197
timestamp 1698431365
transform 1 0 23408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_229
timestamp 1698431365
transform 1 0 26992 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_239
timestamp 1698431365
transform 1 0 28112 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_241
timestamp 1698431365
transform 1 0 28336 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_300
timestamp 1698431365
transform 1 0 34944 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_316
timestamp 1698431365
transform 1 0 36736 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_324
timestamp 1698431365
transform 1 0 37632 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_328
timestamp 1698431365
transform 1 0 38080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_330
timestamp 1698431365
transform 1 0 38304 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_333
timestamp 1698431365
transform 1 0 38640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_10
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_14
timestamp 1698431365
transform 1 0 2912 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_30
timestamp 1698431365
transform 1 0 4704 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_45
timestamp 1698431365
transform 1 0 6384 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_49
timestamp 1698431365
transform 1 0 6832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_66
timestamp 1698431365
transform 1 0 8736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_68
timestamp 1698431365
transform 1 0 8960 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_103
timestamp 1698431365
transform 1 0 12880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_113
timestamp 1698431365
transform 1 0 14000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_153
timestamp 1698431365
transform 1 0 18480 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_157
timestamp 1698431365
transform 1 0 18928 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_249
timestamp 1698431365
transform 1 0 29232 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_302
timestamp 1698431365
transform 1 0 35168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_306
timestamp 1698431365
transform 1 0 35616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_310
timestamp 1698431365
transform 1 0 36064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_333
timestamp 1698431365
transform 1 0 38640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_8
timestamp 1698431365
transform 1 0 2240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_12
timestamp 1698431365
transform 1 0 2688 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_47
timestamp 1698431365
transform 1 0 6608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_51
timestamp 1698431365
transform 1 0 7056 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_55
timestamp 1698431365
transform 1 0 7504 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_57
timestamp 1698431365
transform 1 0 7728 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698431365
transform 1 0 10752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_86
timestamp 1698431365
transform 1 0 10976 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_127
timestamp 1698431365
transform 1 0 15568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_131
timestamp 1698431365
transform 1 0 16016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_133
timestamp 1698431365
transform 1 0 16240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_151
timestamp 1698431365
transform 1 0 18256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_166
timestamp 1698431365
transform 1 0 19936 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_214
timestamp 1698431365
transform 1 0 25312 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_300
timestamp 1698431365
transform 1 0 34944 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_302
timestamp 1698431365
transform 1 0 35168 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_318
timestamp 1698431365
transform 1 0 36960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_322
timestamp 1698431365
transform 1 0 37408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_338
timestamp 1698431365
transform 1 0 39200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698431365
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698431365
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_16
timestamp 1698431365
transform 1 0 3136 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_24
timestamp 1698431365
transform 1 0 4032 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_50
timestamp 1698431365
transform 1 0 6944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_69
timestamp 1698431365
transform 1 0 9072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_76
timestamp 1698431365
transform 1 0 9856 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_122
timestamp 1698431365
transform 1 0 15008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_126
timestamp 1698431365
transform 1 0 15456 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_130
timestamp 1698431365
transform 1 0 15904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_170
timestamp 1698431365
transform 1 0 20384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_183
timestamp 1698431365
transform 1 0 21840 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_198
timestamp 1698431365
transform 1 0 23520 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_202
timestamp 1698431365
transform 1 0 23968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_206
timestamp 1698431365
transform 1 0 24416 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_249
timestamp 1698431365
transform 1 0 29232 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_333
timestamp 1698431365
transform 1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_345
timestamp 1698431365
transform 1 0 39984 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_16
timestamp 1698431365
transform 1 0 3136 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_32
timestamp 1698431365
transform 1 0 4928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_40
timestamp 1698431365
transform 1 0 5824 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_44
timestamp 1698431365
transform 1 0 6272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_47
timestamp 1698431365
transform 1 0 6608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_49
timestamp 1698431365
transform 1 0 6832 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_52
timestamp 1698431365
transform 1 0 7168 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_76
timestamp 1698431365
transform 1 0 9856 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_128
timestamp 1698431365
transform 1 0 15680 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_133
timestamp 1698431365
transform 1 0 16240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_137
timestamp 1698431365
transform 1 0 16688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698431365
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_156
timestamp 1698431365
transform 1 0 18816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_158
timestamp 1698431365
transform 1 0 19040 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_163
timestamp 1698431365
transform 1 0 19600 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_167
timestamp 1698431365
transform 1 0 20048 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_175
timestamp 1698431365
transform 1 0 20944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_177
timestamp 1698431365
transform 1 0 21168 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_203
timestamp 1698431365
transform 1 0 24080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_220
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_222
timestamp 1698431365
transform 1 0 26208 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_239
timestamp 1698431365
transform 1 0 28112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_243
timestamp 1698431365
transform 1 0 28560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_255
timestamp 1698431365
transform 1 0 29904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_257
timestamp 1698431365
transform 1 0 30128 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_264
timestamp 1698431365
transform 1 0 30912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_268
timestamp 1698431365
transform 1 0 31360 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_293
timestamp 1698431365
transform 1 0 34160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_297
timestamp 1698431365
transform 1 0 34608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_301
timestamp 1698431365
transform 1 0 35056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_305
timestamp 1698431365
transform 1 0 35504 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_321
timestamp 1698431365
transform 1 0 37296 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_329
timestamp 1698431365
transform 1 0 38192 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_333
timestamp 1698431365
transform 1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_53
timestamp 1698431365
transform 1 0 7280 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_56
timestamp 1698431365
transform 1 0 7616 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_60
timestamp 1698431365
transform 1 0 8064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_62
timestamp 1698431365
transform 1 0 8288 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_65
timestamp 1698431365
transform 1 0 8624 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_73
timestamp 1698431365
transform 1 0 9520 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_77
timestamp 1698431365
transform 1 0 9968 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_92
timestamp 1698431365
transform 1 0 11648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_94
timestamp 1698431365
transform 1 0 11872 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_103
timestamp 1698431365
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_155
timestamp 1698431365
transform 1 0 18704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_159
timestamp 1698431365
transform 1 0 19152 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_163
timestamp 1698431365
transform 1 0 19600 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_213
timestamp 1698431365
transform 1 0 25200 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_217
timestamp 1698431365
transform 1 0 25648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_231
timestamp 1698431365
transform 1 0 27216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_262
timestamp 1698431365
transform 1 0 30688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_266
timestamp 1698431365
transform 1 0 31136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_280
timestamp 1698431365
transform 1 0 32704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_284
timestamp 1698431365
transform 1 0 33152 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_288
timestamp 1698431365
transform 1 0 33600 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_292
timestamp 1698431365
transform 1 0 34048 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_296
timestamp 1698431365
transform 1 0 34496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_300
timestamp 1698431365
transform 1 0 34944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_304
timestamp 1698431365
transform 1 0 35392 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_18
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_58
timestamp 1698431365
transform 1 0 7840 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_62
timestamp 1698431365
transform 1 0 8288 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_76
timestamp 1698431365
transform 1 0 9856 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_86
timestamp 1698431365
transform 1 0 10976 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_128
timestamp 1698431365
transform 1 0 15680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_132
timestamp 1698431365
transform 1 0 16128 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698431365
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_148
timestamp 1698431365
transform 1 0 17920 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_203
timestamp 1698431365
transform 1 0 24080 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698431365
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_216
timestamp 1698431365
transform 1 0 25536 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_220
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_222
timestamp 1698431365
transform 1 0 26208 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_265
timestamp 1698431365
transform 1 0 31024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_267
timestamp 1698431365
transform 1 0 31248 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_287
timestamp 1698431365
transform 1 0 33488 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_323
timestamp 1698431365
transform 1 0 37520 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_339
timestamp 1698431365
transform 1 0 39312 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_347
timestamp 1698431365
transform 1 0 40208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_16
timestamp 1698431365
transform 1 0 3136 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_32
timestamp 1698431365
transform 1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_88
timestamp 1698431365
transform 1 0 11200 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_92
timestamp 1698431365
transform 1 0 11648 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_96
timestamp 1698431365
transform 1 0 12096 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_98
timestamp 1698431365
transform 1 0 12320 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_116
timestamp 1698431365
transform 1 0 14336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_120
timestamp 1698431365
transform 1 0 14784 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_150
timestamp 1698431365
transform 1 0 18144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_154
timestamp 1698431365
transform 1 0 18592 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_160
timestamp 1698431365
transform 1 0 19264 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_164
timestamp 1698431365
transform 1 0 19712 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_168
timestamp 1698431365
transform 1 0 20160 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698431365
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_189
timestamp 1698431365
transform 1 0 22512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_192
timestamp 1698431365
transform 1 0 22848 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_227
timestamp 1698431365
transform 1 0 26768 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_257
timestamp 1698431365
transform 1 0 30128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_261
timestamp 1698431365
transform 1 0 30576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_263
timestamp 1698431365
transform 1 0 30800 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_281
timestamp 1698431365
transform 1 0 32816 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_321
timestamp 1698431365
transform 1 0 37296 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_325
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_8
timestamp 1698431365
transform 1 0 2240 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_12
timestamp 1698431365
transform 1 0 2688 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_28
timestamp 1698431365
transform 1 0 4480 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_32
timestamp 1698431365
transform 1 0 4928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_34
timestamp 1698431365
transform 1 0 5152 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_45
timestamp 1698431365
transform 1 0 6384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_49
timestamp 1698431365
transform 1 0 6832 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_88
timestamp 1698431365
transform 1 0 11200 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_104
timestamp 1698431365
transform 1 0 12992 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_121
timestamp 1698431365
transform 1 0 14896 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_137
timestamp 1698431365
transform 1 0 16688 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698431365
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_173
timestamp 1698431365
transform 1 0 20720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_177
timestamp 1698431365
transform 1 0 21168 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_193
timestamp 1698431365
transform 1 0 22960 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_201
timestamp 1698431365
transform 1 0 23856 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_203
timestamp 1698431365
transform 1 0 24080 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_216
timestamp 1698431365
transform 1 0 25536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_272
timestamp 1698431365
transform 1 0 31808 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_306
timestamp 1698431365
transform 1 0 35616 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_310
timestamp 1698431365
transform 1 0 36064 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_326
timestamp 1698431365
transform 1 0 37856 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_334
timestamp 1698431365
transform 1 0 38752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_16
timestamp 1698431365
transform 1 0 3136 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_32
timestamp 1698431365
transform 1 0 4928 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_84
timestamp 1698431365
transform 1 0 10752 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_92
timestamp 1698431365
transform 1 0 11648 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_103
timestamp 1698431365
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_109
timestamp 1698431365
transform 1 0 13552 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_183
timestamp 1698431365
transform 1 0 21840 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_187
timestamp 1698431365
transform 1 0 22288 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_207
timestamp 1698431365
transform 1 0 24528 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_209
timestamp 1698431365
transform 1 0 24752 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_212
timestamp 1698431365
transform 1 0 25088 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_243
timestamp 1698431365
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_251
timestamp 1698431365
transform 1 0 29456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_253
timestamp 1698431365
transform 1 0 29680 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_256
timestamp 1698431365
transform 1 0 30016 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_268
timestamp 1698431365
transform 1 0 31360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_270
timestamp 1698431365
transform 1 0 31584 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_308
timestamp 1698431365
transform 1 0 35840 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_312
timestamp 1698431365
transform 1 0 36288 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_49
timestamp 1698431365
transform 1 0 6832 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_93
timestamp 1698431365
transform 1 0 11760 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_129
timestamp 1698431365
transform 1 0 15792 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_133
timestamp 1698431365
transform 1 0 16240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_177
timestamp 1698431365
transform 1 0 21168 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_185
timestamp 1698431365
transform 1 0 22064 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_201
timestamp 1698431365
transform 1 0 23856 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_216
timestamp 1698431365
transform 1 0 25536 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_218
timestamp 1698431365
transform 1 0 25760 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_247
timestamp 1698431365
transform 1 0 29008 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_255
timestamp 1698431365
transform 1 0 29904 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_259
timestamp 1698431365
transform 1 0 30352 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_261
timestamp 1698431365
transform 1 0 30576 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_264
timestamp 1698431365
transform 1 0 30912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_290
timestamp 1698431365
transform 1 0 33824 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_322
timestamp 1698431365
transform 1 0 37408 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_338
timestamp 1698431365
transform 1 0 39200 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_342
timestamp 1698431365
transform 1 0 39648 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_345
timestamp 1698431365
transform 1 0 39984 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_8
timestamp 1698431365
transform 1 0 2240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_12
timestamp 1698431365
transform 1 0 2688 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_28
timestamp 1698431365
transform 1 0 4480 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_32
timestamp 1698431365
transform 1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_42
timestamp 1698431365
transform 1 0 6048 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_46
timestamp 1698431365
transform 1 0 6496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_48
timestamp 1698431365
transform 1 0 6720 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_51
timestamp 1698431365
transform 1 0 7056 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_62
timestamp 1698431365
transform 1 0 8288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_74
timestamp 1698431365
transform 1 0 9632 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_82
timestamp 1698431365
transform 1 0 10528 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_86
timestamp 1698431365
transform 1 0 10976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_88
timestamp 1698431365
transform 1 0 11200 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_94
timestamp 1698431365
transform 1 0 11872 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_102
timestamp 1698431365
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_147
timestamp 1698431365
transform 1 0 17808 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_149
timestamp 1698431365
transform 1 0 18032 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_158
timestamp 1698431365
transform 1 0 19040 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_163
timestamp 1698431365
transform 1 0 19600 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_181
timestamp 1698431365
transform 1 0 21616 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_183
timestamp 1698431365
transform 1 0 21840 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_208
timestamp 1698431365
transform 1 0 24640 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_216
timestamp 1698431365
transform 1 0 25536 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_232
timestamp 1698431365
transform 1 0 27328 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_256
timestamp 1698431365
transform 1 0 30016 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_293
timestamp 1698431365
transform 1 0 34160 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_309
timestamp 1698431365
transform 1 0 35952 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_313
timestamp 1698431365
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_333
timestamp 1698431365
transform 1 0 38640 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_34
timestamp 1698431365
transform 1 0 5152 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_44
timestamp 1698431365
transform 1 0 6272 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_48
timestamp 1698431365
transform 1 0 6720 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_51
timestamp 1698431365
transform 1 0 7056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_67
timestamp 1698431365
transform 1 0 8848 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_74
timestamp 1698431365
transform 1 0 9632 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_88
timestamp 1698431365
transform 1 0 11200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_92
timestamp 1698431365
transform 1 0 11648 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_96
timestamp 1698431365
transform 1 0 12096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_98
timestamp 1698431365
transform 1 0 12320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_116
timestamp 1698431365
transform 1 0 14336 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_126
timestamp 1698431365
transform 1 0 15456 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_144
timestamp 1698431365
transform 1 0 17472 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_177
timestamp 1698431365
transform 1 0 21168 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_185
timestamp 1698431365
transform 1 0 22064 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_193
timestamp 1698431365
transform 1 0 22960 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_199
timestamp 1698431365
transform 1 0 23632 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_209
timestamp 1698431365
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_224
timestamp 1698431365
transform 1 0 26432 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_226
timestamp 1698431365
transform 1 0 26656 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_240
timestamp 1698431365
transform 1 0 28224 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_256
timestamp 1698431365
transform 1 0 30016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_258
timestamp 1698431365
transform 1 0 30240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_295
timestamp 1698431365
transform 1 0 34384 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_327
timestamp 1698431365
transform 1 0 37968 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_343
timestamp 1698431365
transform 1 0 39760 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_347
timestamp 1698431365
transform 1 0 40208 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_53
timestamp 1698431365
transform 1 0 7280 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_99
timestamp 1698431365
transform 1 0 12432 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_103
timestamp 1698431365
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_115
timestamp 1698431365
transform 1 0 14224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_141
timestamp 1698431365
transform 1 0 17136 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_163
timestamp 1698431365
transform 1 0 19600 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_167
timestamp 1698431365
transform 1 0 20048 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_214
timestamp 1698431365
transform 1 0 25312 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_218
timestamp 1698431365
transform 1 0 25760 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_242
timestamp 1698431365
transform 1 0 28448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_244
timestamp 1698431365
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_255
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_257
timestamp 1698431365
transform 1 0 30128 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_305
timestamp 1698431365
transform 1 0 35504 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_18
timestamp 1698431365
transform 1 0 3360 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_20
timestamp 1698431365
transform 1 0 3584 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_55
timestamp 1698431365
transform 1 0 7504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_57
timestamp 1698431365
transform 1 0 7728 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_74
timestamp 1698431365
transform 1 0 9632 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_108
timestamp 1698431365
transform 1 0 13440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_160
timestamp 1698431365
transform 1 0 19264 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_164
timestamp 1698431365
transform 1 0 19712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_248
timestamp 1698431365
transform 1 0 29120 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_252
timestamp 1698431365
transform 1 0 29568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_256
timestamp 1698431365
transform 1 0 30016 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_294
timestamp 1698431365
transform 1 0 34272 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_326
timestamp 1698431365
transform 1 0 37856 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_342
timestamp 1698431365
transform 1 0 39648 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698431365
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698431365
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_45
timestamp 1698431365
transform 1 0 6384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_47
timestamp 1698431365
transform 1 0 6608 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_53
timestamp 1698431365
transform 1 0 7280 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_57
timestamp 1698431365
transform 1 0 7728 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_61
timestamp 1698431365
transform 1 0 8176 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_63
timestamp 1698431365
transform 1 0 8400 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_97
timestamp 1698431365
transform 1 0 12208 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_109
timestamp 1698431365
transform 1 0 13552 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_159
timestamp 1698431365
transform 1 0 19152 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_163
timestamp 1698431365
transform 1 0 19600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_167
timestamp 1698431365
transform 1 0 20048 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_179
timestamp 1698431365
transform 1 0 21392 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_211
timestamp 1698431365
transform 1 0 24976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_215
timestamp 1698431365
transform 1 0 25424 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_219
timestamp 1698431365
transform 1 0 25872 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_223
timestamp 1698431365
transform 1 0 26320 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_236
timestamp 1698431365
transform 1 0 27776 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_242
timestamp 1698431365
transform 1 0 28448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698431365
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_251
timestamp 1698431365
transform 1 0 29456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_255
timestamp 1698431365
transform 1 0 29904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_257
timestamp 1698431365
transform 1 0 30128 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_260
timestamp 1698431365
transform 1 0 30464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_262
timestamp 1698431365
transform 1 0 30688 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_265
timestamp 1698431365
transform 1 0 31024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_284
timestamp 1698431365
transform 1 0 33152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_289
timestamp 1698431365
transform 1 0 33712 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_293
timestamp 1698431365
transform 1 0 34160 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_297
timestamp 1698431365
transform 1 0 34608 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_313
timestamp 1698431365
transform 1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_76
timestamp 1698431365
transform 1 0 9856 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_79
timestamp 1698431365
transform 1 0 10192 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_83
timestamp 1698431365
transform 1 0 10640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_100
timestamp 1698431365
transform 1 0 12544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_104
timestamp 1698431365
transform 1 0 12992 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_107
timestamp 1698431365
transform 1 0 13328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_166
timestamp 1698431365
transform 1 0 19936 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_168
timestamp 1698431365
transform 1 0 20160 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_171
timestamp 1698431365
transform 1 0 20496 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_194
timestamp 1698431365
transform 1 0 23072 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_196
timestamp 1698431365
transform 1 0 23296 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_202
timestamp 1698431365
transform 1 0 23968 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_220
timestamp 1698431365
transform 1 0 25984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_228
timestamp 1698431365
transform 1 0 26880 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_235
timestamp 1698431365
transform 1 0 27664 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_239
timestamp 1698431365
transform 1 0 28112 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_243
timestamp 1698431365
transform 1 0 28560 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_248
timestamp 1698431365
transform 1 0 29120 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_252
timestamp 1698431365
transform 1 0 29568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_256
timestamp 1698431365
transform 1 0 30016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_268
timestamp 1698431365
transform 1 0 31360 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_270
timestamp 1698431365
transform 1 0 31584 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_287
timestamp 1698431365
transform 1 0 33488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_291
timestamp 1698431365
transform 1 0 33936 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_297
timestamp 1698431365
transform 1 0 34608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_301
timestamp 1698431365
transform 1 0 35056 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_333
timestamp 1698431365
transform 1 0 38640 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_53
timestamp 1698431365
transform 1 0 7280 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_61
timestamp 1698431365
transform 1 0 8176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_65
timestamp 1698431365
transform 1 0 8624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_113
timestamp 1698431365
transform 1 0 14000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_115
timestamp 1698431365
transform 1 0 14224 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698431365
transform 1 0 20720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_195
timestamp 1698431365
transform 1 0 23184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_197
timestamp 1698431365
transform 1 0 23408 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_81
timestamp 1698431365
transform 1 0 10416 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_83
timestamp 1698431365
transform 1 0 10640 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_86
timestamp 1698431365
transform 1 0 10976 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_152
timestamp 1698431365
transform 1 0 18368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_217
timestamp 1698431365
transform 1 0 25648 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_261
timestamp 1698431365
transform 1 0 30576 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_286
timestamp 1698431365
transform 1 0 33376 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_290
timestamp 1698431365
transform 1 0 33824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_294
timestamp 1698431365
transform 1 0 34272 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_298
timestamp 1698431365
transform 1 0 34720 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_302
timestamp 1698431365
transform 1 0 35168 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_334
timestamp 1698431365
transform 1 0 38752 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_342
timestamp 1698431365
transform 1 0 39648 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698431365
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698431365
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698431365
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_80
timestamp 1698431365
transform 1 0 10304 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_84
timestamp 1698431365
transform 1 0 10752 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_87
timestamp 1698431365
transform 1 0 11088 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_97
timestamp 1698431365
transform 1 0 12208 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_99
timestamp 1698431365
transform 1 0 12432 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_114
timestamp 1698431365
transform 1 0 14112 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_118
timestamp 1698431365
transform 1 0 14560 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_121
timestamp 1698431365
transform 1 0 14896 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_135
timestamp 1698431365
transform 1 0 16464 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_138
timestamp 1698431365
transform 1 0 16800 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_152
timestamp 1698431365
transform 1 0 18368 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_156
timestamp 1698431365
transform 1 0 18816 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698431365
transform 1 0 20608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698431365
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_189
timestamp 1698431365
transform 1 0 22512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_200
timestamp 1698431365
transform 1 0 23744 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_234
timestamp 1698431365
transform 1 0 27552 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_250
timestamp 1698431365
transform 1 0 29344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_264
timestamp 1698431365
transform 1 0 30912 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_268
timestamp 1698431365
transform 1 0 31360 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_274
timestamp 1698431365
transform 1 0 32032 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_276
timestamp 1698431365
transform 1 0 32256 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_291
timestamp 1698431365
transform 1 0 33936 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698431365
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698431365
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698431365
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698431365
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13888 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input1
timestamp 1698431365
transform -1 0 40432 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input3
timestamp 1698431365
transform 1 0 3136 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input4
timestamp 1698431365
transform 1 0 3136 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input5
timestamp 1698431365
transform 1 0 2464 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input6
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input7
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input10
timestamp 1698431365
transform 1 0 9520 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input11
timestamp 1698431365
transform 1 0 11536 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input12
timestamp 1698431365
transform -1 0 40432 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input13
timestamp 1698431365
transform -1 0 17024 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input14
timestamp 1698431365
transform -1 0 16128 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input15
timestamp 1698431365
transform -1 0 19488 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input16
timestamp 1698431365
transform 1 0 18816 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input17
timestamp 1698431365
transform -1 0 24192 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input18
timestamp 1698431365
transform -1 0 24864 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 27664 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input20
timestamp 1698431365
transform -1 0 30576 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input21
timestamp 1698431365
transform -1 0 32592 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input22
timestamp 1698431365
transform -1 0 39760 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform -1 0 40432 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input24
timestamp 1698431365
transform -1 0 40432 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 40432 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform -1 0 40432 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input27
timestamp 1698431365
transform -1 0 26320 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input28
timestamp 1698431365
transform -1 0 39760 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input29
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 40432 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input31
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input32
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 23856 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output34
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output35 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38864 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output36
timestamp 1698431365
transform 1 0 38864 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output37
timestamp 1698431365
transform 1 0 38864 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output38
timestamp 1698431365
transform 1 0 26320 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output39
timestamp 1698431365
transform 1 0 38864 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output40
timestamp 1698431365
transform 1 0 38864 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output41
timestamp 1698431365
transform -1 0 3136 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output42
timestamp 1698431365
transform -1 0 3136 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output43
timestamp 1698431365
transform -1 0 3136 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output44
timestamp 1698431365
transform -1 0 3136 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output45
timestamp 1698431365
transform -1 0 3136 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output46
timestamp 1698431365
transform -1 0 3136 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output47
timestamp 1698431365
transform -1 0 3136 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output48
timestamp 1698431365
transform -1 0 3136 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output49
timestamp 1698431365
transform 1 0 9184 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output50
timestamp 1698431365
transform -1 0 14112 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output51
timestamp 1698431365
transform 1 0 38864 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output52
timestamp 1698431365
transform 1 0 17248 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output53
timestamp 1698431365
transform -1 0 16464 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output54
timestamp 1698431365
transform -1 0 18368 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output55
timestamp 1698431365
transform -1 0 22512 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output56
timestamp 1698431365
transform -1 0 23744 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output57
timestamp 1698431365
transform -1 0 27552 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output58
timestamp 1698431365
transform 1 0 29792 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output59
timestamp 1698431365
transform 1 0 28224 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output60
timestamp 1698431365
transform -1 0 35616 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output61
timestamp 1698431365
transform -1 0 33936 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output62
timestamp 1698431365
transform 1 0 38864 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output63
timestamp 1698431365
transform 1 0 38864 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output64
timestamp 1698431365
transform 1 0 38864 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output65
timestamp 1698431365
transform 1 0 38864 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output66
timestamp 1698431365
transform 1 0 38864 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output67
timestamp 1698431365
transform 1 0 38864 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output68
timestamp 1698431365
transform 1 0 19264 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output69
timestamp 1698431365
transform -1 0 25984 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output70
timestamp 1698431365
transform -1 0 3136 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output71
timestamp 1698431365
transform -1 0 3136 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output72
timestamp 1698431365
transform 1 0 21616 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output73
timestamp 1698431365
transform 1 0 18256 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698431365
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698431365
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698431365
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698431365
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698431365
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698431365
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698431365
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698431365
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698431365
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 clock
port 0 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 logisim_clock_tree_0_out
port 1 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 ram_addr_o[0]
port 2 nsew signal tristate
flabel metal3 s 41200 16128 42000 16240 0 FreeSans 448 0 0 0 ram_addr_o[1]
port 3 nsew signal tristate
flabel metal3 s 41200 15456 42000 15568 0 FreeSans 448 0 0 0 ram_addr_o[2]
port 4 nsew signal tristate
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 ram_addr_o[3]
port 5 nsew signal tristate
flabel metal3 s 41200 14784 42000 14896 0 FreeSans 448 0 0 0 ram_addr_o[4]
port 6 nsew signal tristate
flabel metal3 s 41200 14112 42000 14224 0 FreeSans 448 0 0 0 ram_data_i[0]
port 7 nsew signal input
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 ram_data_i[10]
port 8 nsew signal input
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 ram_data_i[11]
port 9 nsew signal input
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 ram_data_i[12]
port 10 nsew signal input
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 ram_data_i[13]
port 11 nsew signal input
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 ram_data_i[14]
port 12 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 ram_data_i[15]
port 13 nsew signal input
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 ram_data_i[16]
port 14 nsew signal input
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 ram_data_i[17]
port 15 nsew signal input
flabel metal2 s 9408 41200 9520 42000 0 FreeSans 448 90 0 0 ram_data_i[18]
port 16 nsew signal input
flabel metal2 s 11424 41200 11536 42000 0 FreeSans 448 90 0 0 ram_data_i[19]
port 17 nsew signal input
flabel metal3 s 41200 12768 42000 12880 0 FreeSans 448 0 0 0 ram_data_i[1]
port 18 nsew signal input
flabel metal2 s 17472 41200 17584 42000 0 FreeSans 448 90 0 0 ram_data_i[20]
port 19 nsew signal input
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 ram_data_i[21]
port 20 nsew signal input
flabel metal2 s 18144 41200 18256 42000 0 FreeSans 448 90 0 0 ram_data_i[22]
port 21 nsew signal input
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 ram_data_i[23]
port 22 nsew signal input
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 ram_data_i[24]
port 23 nsew signal input
flabel metal2 s 23520 41200 23632 42000 0 FreeSans 448 90 0 0 ram_data_i[25]
port 24 nsew signal input
flabel metal2 s 26880 41200 26992 42000 0 FreeSans 448 90 0 0 ram_data_i[26]
port 25 nsew signal input
flabel metal2 s 27552 41200 27664 42000 0 FreeSans 448 90 0 0 ram_data_i[27]
port 26 nsew signal input
flabel metal2 s 31584 41200 31696 42000 0 FreeSans 448 90 0 0 ram_data_i[28]
port 27 nsew signal input
flabel metal3 s 41200 31584 42000 31696 0 FreeSans 448 0 0 0 ram_data_i[29]
port 28 nsew signal input
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 ram_data_i[2]
port 29 nsew signal input
flabel metal3 s 41200 30912 42000 31024 0 FreeSans 448 0 0 0 ram_data_i[30]
port 30 nsew signal input
flabel metal3 s 41200 28224 42000 28336 0 FreeSans 448 0 0 0 ram_data_i[31]
port 31 nsew signal input
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 ram_data_i[3]
port 32 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 ram_data_i[4]
port 33 nsew signal input
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 ram_data_i[5]
port 34 nsew signal input
flabel metal2 s 21504 41200 21616 42000 0 FreeSans 448 90 0 0 ram_data_i[6]
port 35 nsew signal input
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 ram_data_i[7]
port 36 nsew signal input
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 ram_data_i[8]
port 37 nsew signal input
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 ram_data_i[9]
port 38 nsew signal input
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 ram_data_o[0]
port 39 nsew signal tristate
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 ram_data_o[10]
port 40 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 ram_data_o[11]
port 41 nsew signal tristate
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 ram_data_o[12]
port 42 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 ram_data_o[13]
port 43 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 ram_data_o[14]
port 44 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 ram_data_o[15]
port 45 nsew signal tristate
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 ram_data_o[16]
port 46 nsew signal tristate
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 ram_data_o[17]
port 47 nsew signal tristate
flabel metal2 s 8736 41200 8848 42000 0 FreeSans 448 90 0 0 ram_data_o[18]
port 48 nsew signal tristate
flabel metal2 s 12096 41200 12208 42000 0 FreeSans 448 90 0 0 ram_data_o[19]
port 49 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 ram_data_o[1]
port 50 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 ram_data_o[20]
port 51 nsew signal tristate
flabel metal2 s 14784 41200 14896 42000 0 FreeSans 448 90 0 0 ram_data_o[21]
port 52 nsew signal tristate
flabel metal2 s 16128 41200 16240 42000 0 FreeSans 448 90 0 0 ram_data_o[22]
port 53 nsew signal tristate
flabel metal2 s 20832 41200 20944 42000 0 FreeSans 448 90 0 0 ram_data_o[23]
port 54 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 ram_data_o[24]
port 55 nsew signal tristate
flabel metal2 s 25536 41200 25648 42000 0 FreeSans 448 90 0 0 ram_data_o[25]
port 56 nsew signal tristate
flabel metal2 s 28896 41200 29008 42000 0 FreeSans 448 90 0 0 ram_data_o[26]
port 57 nsew signal tristate
flabel metal2 s 26208 41200 26320 42000 0 FreeSans 448 90 0 0 ram_data_o[27]
port 58 nsew signal tristate
flabel metal2 s 34272 41200 34384 42000 0 FreeSans 448 90 0 0 ram_data_o[28]
port 59 nsew signal tristate
flabel metal2 s 32256 41200 32368 42000 0 FreeSans 448 90 0 0 ram_data_o[29]
port 60 nsew signal tristate
flabel metal3 s 41200 25536 42000 25648 0 FreeSans 448 0 0 0 ram_data_o[2]
port 61 nsew signal tristate
flabel metal3 s 41200 28896 42000 29008 0 FreeSans 448 0 0 0 ram_data_o[30]
port 62 nsew signal tristate
flabel metal3 s 41200 13440 42000 13552 0 FreeSans 448 0 0 0 ram_data_o[31]
port 63 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 ram_data_o[3]
port 64 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 ram_data_o[4]
port 65 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 ram_data_o[5]
port 66 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 ram_data_o[6]
port 67 nsew signal tristate
flabel metal2 s 24192 41200 24304 42000 0 FreeSans 448 90 0 0 ram_data_o[7]
port 68 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 ram_data_o[8]
port 69 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 ram_data_o[9]
port 70 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 ram_rw_en_o
port 71 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 reset_i
port 72 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 stop_lamp_o
port 73 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 74 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 74 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 75 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 14840 10248 14840 10248 0 _0000_
rlabel metal2 37800 13496 37800 13496 0 _0001_
rlabel metal2 38416 10584 38416 10584 0 _0002_
rlabel metal2 35784 7840 35784 7840 0 _0003_
rlabel metal3 30296 7560 30296 7560 0 _0004_
rlabel metal2 26824 6496 26824 6496 0 _0005_
rlabel metal2 37856 21784 37856 21784 0 _0006_
rlabel metal2 37688 19768 37688 19768 0 _0007_
rlabel metal2 36680 24976 36680 24976 0 _0008_
rlabel metal2 29624 24472 29624 24472 0 _0009_
rlabel metal2 27440 24920 27440 24920 0 _0010_
rlabel metal2 23576 18760 23576 18760 0 _0011_
rlabel metal2 19544 25704 19544 25704 0 _0012_
rlabel metal2 23912 26656 23912 26656 0 _0013_
rlabel metal2 17920 23688 17920 23688 0 _0014_
rlabel metal3 20832 18984 20832 18984 0 _0015_
rlabel metal3 14000 15512 14000 15512 0 _0016_
rlabel metal2 9688 15680 9688 15680 0 _0017_
rlabel metal2 4760 21952 4760 21952 0 _0018_
rlabel metal2 4984 18256 4984 18256 0 _0019_
rlabel metal3 4312 24920 4312 24920 0 _0020_
rlabel metal2 14728 26880 14728 26880 0 _0021_
rlabel metal3 7168 28056 7168 28056 0 _0022_
rlabel metal2 3304 31360 3304 31360 0 _0023_
rlabel metal3 6832 33544 6832 33544 0 _0024_
rlabel metal3 12376 36232 12376 36232 0 _0025_
rlabel metal3 20048 36232 20048 36232 0 _0026_
rlabel metal2 14056 36008 14056 36008 0 _0027_
rlabel metal2 16072 26656 16072 26656 0 _0028_
rlabel metal2 21840 28056 21840 28056 0 _0029_
rlabel metal2 22904 37072 22904 37072 0 _0030_
rlabel metal2 26600 36064 26600 36064 0 _0031_
rlabel metal2 28952 36680 28952 36680 0 _0032_
rlabel metal2 25928 28840 25928 28840 0 _0033_
rlabel metal2 34440 36064 34440 36064 0 _0034_
rlabel metal3 31472 36344 31472 36344 0 _0035_
rlabel metal2 36960 28056 36960 28056 0 _0036_
rlabel metal3 30240 28056 30240 28056 0 _0037_
rlabel metal3 33712 17416 33712 17416 0 _0038_
rlabel metal2 36232 16632 36232 16632 0 _0039_
rlabel metal2 29512 16464 29512 16464 0 _0040_
rlabel metal3 25536 8008 25536 8008 0 _0041_
rlabel metal2 26936 17248 26936 17248 0 _0042_
rlabel metal2 24472 16240 24472 16240 0 _0043_
rlabel metal2 17976 14672 17976 14672 0 _0044_
rlabel metal2 16856 15680 16856 15680 0 _0045_
rlabel metal2 21336 8848 21336 8848 0 _0046_
rlabel metal2 21336 7280 21336 7280 0 _0047_
rlabel metal3 20384 10024 20384 10024 0 _0048_
rlabel metal2 18088 11312 18088 11312 0 _0049_
rlabel metal2 34216 13104 34216 13104 0 _0050_
rlabel metal2 35336 10752 35336 10752 0 _0051_
rlabel metal2 33208 8792 33208 8792 0 _0052_
rlabel metal2 30912 7448 30912 7448 0 _0053_
rlabel metal2 24472 7392 24472 7392 0 _0054_
rlabel metal2 34888 21616 34888 21616 0 _0055_
rlabel metal2 35112 19544 35112 19544 0 _0056_
rlabel metal2 33432 25648 33432 25648 0 _0057_
rlabel metal2 28280 24864 28280 24864 0 _0058_
rlabel metal2 26824 25200 26824 25200 0 _0059_
rlabel metal2 21000 20272 21000 20272 0 _0060_
rlabel metal3 18032 24920 18032 24920 0 _0061_
rlabel metal2 21896 27328 21896 27328 0 _0062_
rlabel metal3 17528 23184 17528 23184 0 _0063_
rlabel metal3 17304 19208 17304 19208 0 _0064_
rlabel metal2 11144 15624 11144 15624 0 _0065_
rlabel metal2 7336 16408 7336 16408 0 _0066_
rlabel metal2 4760 20888 4760 20888 0 _0067_
rlabel metal2 2632 18368 2632 18368 0 _0068_
rlabel metal2 5824 24696 5824 24696 0 _0069_
rlabel metal2 12264 27496 12264 27496 0 _0070_
rlabel metal2 4312 28112 4312 28112 0 _0071_
rlabel metal2 5712 29624 5712 29624 0 _0072_
rlabel metal3 5264 33432 5264 33432 0 _0073_
rlabel metal3 10472 35896 10472 35896 0 _0074_
rlabel metal2 16408 35840 16408 35840 0 _0075_
rlabel metal2 13496 36512 13496 36512 0 _0076_
rlabel metal2 14056 26208 14056 26208 0 _0077_
rlabel metal2 19544 28616 19544 28616 0 _0078_
rlabel metal2 21448 36904 21448 36904 0 _0079_
rlabel metal2 25368 36176 25368 36176 0 _0080_
rlabel metal2 26600 36904 26600 36904 0 _0081_
rlabel metal2 23688 29064 23688 29064 0 _0082_
rlabel metal2 32032 35896 32032 35896 0 _0083_
rlabel metal2 30744 36176 30744 36176 0 _0084_
rlabel metal2 34440 28112 34440 28112 0 _0085_
rlabel metal2 27272 27944 27272 27944 0 _0086_
rlabel metal2 31192 16912 31192 16912 0 _0087_
rlabel metal2 34104 16968 34104 16968 0 _0088_
rlabel metal2 27328 15288 27328 15288 0 _0089_
rlabel metal3 23072 7560 23072 7560 0 _0090_
rlabel metal3 25256 15512 25256 15512 0 _0091_
rlabel metal2 21560 14504 21560 14504 0 _0092_
rlabel metal2 15736 15148 15736 15148 0 _0093_
rlabel metal2 15176 16240 15176 16240 0 _0094_
rlabel metal2 12824 11424 12824 11424 0 _0095_
rlabel metal3 17080 13048 17080 13048 0 _0096_
rlabel metal2 10360 10920 10360 10920 0 _0097_
rlabel metal2 5992 11816 5992 11816 0 _0098_
rlabel metal2 2968 13440 2968 13440 0 _0099_
rlabel metal2 8232 14056 8232 14056 0 _0100_
rlabel metal2 21000 11816 21000 11816 0 _0101_
rlabel metal2 21112 16128 21112 16128 0 _0102_
rlabel metal2 26264 13440 26264 13440 0 _0103_
rlabel metal2 19264 12936 19264 12936 0 _0104_
rlabel metal2 18312 12600 18312 12600 0 _0105_
rlabel metal2 15176 21672 15176 21672 0 _0106_
rlabel metal2 23128 10925 23128 10925 0 _0107_
rlabel metal3 21728 18312 21728 18312 0 _0108_
rlabel metal3 15792 16744 15792 16744 0 _0109_
rlabel metal3 16632 16856 16632 16856 0 _0110_
rlabel metal2 15848 16016 15848 16016 0 _0111_
rlabel metal3 16800 15288 16800 15288 0 _0112_
rlabel metal2 21672 14056 21672 14056 0 _0113_
rlabel metal2 21896 16632 21896 16632 0 _0114_
rlabel metal2 25928 16128 25928 16128 0 _0115_
rlabel metal2 26376 15568 26376 15568 0 _0116_
rlabel metal2 28280 23856 28280 23856 0 _0117_
rlabel metal3 24584 7560 24584 7560 0 _0118_
rlabel metal2 30520 15960 30520 15960 0 _0119_
rlabel metal2 28168 15904 28168 15904 0 _0120_
rlabel metal2 33880 19320 33880 19320 0 _0121_
rlabel metal2 34328 16856 34328 16856 0 _0122_
rlabel metal2 32760 18592 32760 18592 0 _0123_
rlabel metal2 31752 16352 31752 16352 0 _0124_
rlabel metal2 19656 16352 19656 16352 0 _0125_
rlabel metal2 26376 22064 26376 22064 0 _0126_
rlabel metal2 33320 28448 33320 28448 0 _0127_
rlabel metal3 31976 28056 31976 28056 0 _0128_
rlabel metal2 19208 30632 19208 30632 0 _0129_
rlabel metal2 21448 30632 21448 30632 0 _0130_
rlabel metal2 17752 29624 17752 29624 0 _0131_
rlabel metal2 18032 30968 18032 30968 0 _0132_
rlabel metal3 15848 34664 15848 34664 0 _0133_
rlabel metal2 13944 34160 13944 34160 0 _0134_
rlabel metal2 14504 35672 14504 35672 0 _0135_
rlabel metal2 14616 33656 14616 33656 0 _0136_
rlabel metal2 14952 32200 14952 32200 0 _0137_
rlabel metal2 9352 33992 9352 33992 0 _0138_
rlabel metal3 13384 31640 13384 31640 0 _0139_
rlabel metal2 18424 32928 18424 32928 0 _0140_
rlabel metal2 13608 31808 13608 31808 0 _0141_
rlabel metal2 10136 32592 10136 32592 0 _0142_
rlabel metal2 10808 34048 10808 34048 0 _0143_
rlabel metal3 11872 31640 11872 31640 0 _0144_
rlabel metal3 8008 31080 8008 31080 0 _0145_
rlabel metal2 9464 30800 9464 30800 0 _0146_
rlabel metal2 8792 31416 8792 31416 0 _0147_
rlabel metal2 9352 29904 9352 29904 0 _0148_
rlabel metal2 8904 30520 8904 30520 0 _0149_
rlabel metal2 11480 30632 11480 30632 0 _0150_
rlabel metal2 13608 32200 13608 32200 0 _0151_
rlabel metal3 13776 31080 13776 31080 0 _0152_
rlabel metal2 14728 32256 14728 32256 0 _0153_
rlabel metal2 15624 34496 15624 34496 0 _0154_
rlabel metal3 17696 35784 17696 35784 0 _0155_
rlabel metal2 14952 34720 14952 34720 0 _0156_
rlabel metal3 18648 34608 18648 34608 0 _0157_
rlabel metal2 15176 32816 15176 32816 0 _0158_
rlabel metal2 14840 31752 14840 31752 0 _0159_
rlabel metal3 18592 30968 18592 30968 0 _0160_
rlabel metal2 20664 31136 20664 31136 0 _0161_
rlabel metal3 21616 31752 21616 31752 0 _0162_
rlabel metal2 11144 23520 11144 23520 0 _0163_
rlabel metal2 8008 25312 8008 25312 0 _0164_
rlabel metal3 11088 23912 11088 23912 0 _0165_
rlabel metal2 7336 23184 7336 23184 0 _0166_
rlabel metal2 8344 23184 8344 23184 0 _0167_
rlabel metal2 11480 22736 11480 22736 0 _0168_
rlabel metal2 10808 18928 10808 18928 0 _0169_
rlabel metal2 12824 18704 12824 18704 0 _0170_
rlabel metal2 11536 17752 11536 17752 0 _0171_
rlabel metal2 12152 19992 12152 19992 0 _0172_
rlabel metal3 15792 18424 15792 18424 0 _0173_
rlabel metal2 15960 21280 15960 21280 0 _0174_
rlabel metal2 16464 20776 16464 20776 0 _0175_
rlabel metal2 15400 18872 15400 18872 0 _0176_
rlabel metal2 13944 20048 13944 20048 0 _0177_
rlabel metal2 12152 17528 12152 17528 0 _0178_
rlabel metal2 12600 16800 12600 16800 0 _0179_
rlabel metal2 11928 18480 11928 18480 0 _0180_
rlabel metal2 11648 20664 11648 20664 0 _0181_
rlabel metal2 12376 21280 12376 21280 0 _0182_
rlabel metal2 22120 25088 22120 25088 0 _0183_
rlabel metal2 23352 25256 23352 25256 0 _0184_
rlabel metal2 20272 24024 20272 24024 0 _0185_
rlabel metal3 23520 23800 23520 23800 0 _0186_
rlabel metal2 24472 23408 24472 23408 0 _0187_
rlabel metal2 25704 22792 25704 22792 0 _0188_
rlabel metal3 29400 23912 29400 23912 0 _0189_
rlabel metal3 29344 22456 29344 22456 0 _0190_
rlabel metal2 33544 24192 33544 24192 0 _0191_
rlabel metal2 31192 23352 31192 23352 0 _0192_
rlabel metal3 34384 23240 34384 23240 0 _0193_
rlabel metal2 34440 20496 34440 20496 0 _0194_
rlabel metal2 34048 22232 34048 22232 0 _0195_
rlabel metal2 34216 24584 34216 24584 0 _0196_
rlabel metal2 31752 25032 31752 25032 0 _0197_
rlabel metal2 33208 23800 33208 23800 0 _0198_
rlabel metal2 32200 23240 32200 23240 0 _0199_
rlabel metal3 28896 21672 28896 21672 0 _0200_
rlabel metal2 28616 22848 28616 22848 0 _0201_
rlabel metal2 26824 23072 26824 23072 0 _0202_
rlabel metal2 23016 23576 23016 23576 0 _0203_
rlabel metal3 24864 19432 24864 19432 0 _0204_
rlabel metal3 25564 21336 25564 21336 0 _0205_
rlabel metal2 26600 22456 26600 22456 0 _0206_
rlabel metal2 25704 20496 25704 20496 0 _0207_
rlabel metal2 21672 22848 21672 22848 0 _0208_
rlabel metal2 23408 24696 23408 24696 0 _0209_
rlabel metal2 21560 25032 21560 25032 0 _0210_
rlabel metal2 23240 24248 23240 24248 0 _0211_
rlabel metal2 23352 23016 23352 23016 0 _0212_
rlabel metal2 15960 22400 15960 22400 0 _0213_
rlabel metal2 15400 20328 15400 20328 0 _0214_
rlabel metal2 16184 22792 16184 22792 0 _0215_
rlabel metal2 13496 21056 13496 21056 0 _0216_
rlabel metal2 12712 21672 12712 21672 0 _0217_
rlabel metal3 12208 22120 12208 22120 0 _0218_
rlabel metal3 13496 21784 13496 21784 0 _0219_
rlabel metal2 10696 24416 10696 24416 0 _0220_
rlabel metal2 6160 18648 6160 18648 0 _0221_
rlabel metal2 5768 20272 5768 20272 0 _0222_
rlabel metal2 6216 20272 6216 20272 0 _0223_
rlabel metal3 6720 20776 6720 20776 0 _0224_
rlabel metal2 6888 18200 6888 18200 0 _0225_
rlabel metal2 8792 22736 8792 22736 0 _0226_
rlabel metal2 10024 23520 10024 23520 0 _0227_
rlabel metal2 12712 25984 12712 25984 0 _0228_
rlabel metal2 9576 25872 9576 25872 0 _0229_
rlabel metal3 12096 26488 12096 26488 0 _0230_
rlabel metal2 13608 28336 13608 28336 0 _0231_
rlabel metal2 8400 29512 8400 29512 0 _0232_
rlabel metal3 9240 28728 9240 28728 0 _0233_
rlabel metal2 10920 29848 10920 29848 0 _0234_
rlabel metal2 10472 30240 10472 30240 0 _0235_
rlabel metal2 14056 30240 14056 30240 0 _0236_
rlabel metal2 18648 30296 18648 30296 0 _0237_
rlabel metal2 15512 29848 15512 29848 0 _0238_
rlabel metal2 14728 29680 14728 29680 0 _0239_
rlabel metal2 22232 30912 22232 30912 0 _0240_
rlabel metal2 29288 30520 29288 30520 0 _0241_
rlabel metal2 25928 30856 25928 30856 0 _0242_
rlabel metal3 26572 34104 26572 34104 0 _0243_
rlabel metal3 26040 31584 26040 31584 0 _0244_
rlabel metal3 26152 31752 26152 31752 0 _0245_
rlabel metal2 24584 35392 24584 35392 0 _0246_
rlabel metal2 23240 33376 23240 33376 0 _0247_
rlabel metal3 23240 34104 23240 34104 0 _0248_
rlabel metal2 23016 32536 23016 32536 0 _0249_
rlabel metal2 23800 32536 23800 32536 0 _0250_
rlabel metal2 23912 31808 23912 31808 0 _0251_
rlabel metal3 23352 31472 23352 31472 0 _0252_
rlabel metal2 26824 31360 26824 31360 0 _0253_
rlabel metal2 27944 32032 27944 32032 0 _0254_
rlabel metal2 26152 33488 26152 33488 0 _0255_
rlabel metal2 27384 32816 27384 32816 0 _0256_
rlabel metal2 25032 34216 25032 34216 0 _0257_
rlabel metal3 21728 35112 21728 35112 0 _0258_
rlabel metal3 24696 34160 24696 34160 0 _0259_
rlabel metal2 25144 33432 25144 33432 0 _0260_
rlabel metal2 24696 32200 24696 32200 0 _0261_
rlabel metal3 27272 31640 27272 31640 0 _0262_
rlabel metal2 30520 32200 30520 32200 0 _0263_
rlabel metal3 33936 32536 33936 32536 0 _0264_
rlabel metal3 31416 33208 31416 33208 0 _0265_
rlabel metal3 34384 34104 34384 34104 0 _0266_
rlabel metal2 33768 33488 33768 33488 0 _0267_
rlabel metal2 31304 32032 31304 32032 0 _0268_
rlabel metal2 32200 31024 32200 31024 0 _0269_
rlabel metal2 33880 32088 33880 32088 0 _0270_
rlabel metal2 32984 33656 32984 33656 0 _0271_
rlabel metal2 33656 31752 33656 31752 0 _0272_
rlabel metal2 33096 31360 33096 31360 0 _0273_
rlabel metal3 34328 30968 34328 30968 0 _0274_
rlabel metal3 32256 30184 32256 30184 0 _0275_
rlabel metal3 31080 27720 31080 27720 0 _0276_
rlabel metal2 31752 27608 31752 27608 0 _0277_
rlabel metal2 31080 29400 31080 29400 0 _0278_
rlabel metal2 19600 15288 19600 15288 0 _0279_
rlabel metal2 20160 15512 20160 15512 0 _0280_
rlabel metal3 25704 17192 25704 17192 0 _0281_
rlabel metal3 28952 31640 28952 31640 0 _0282_
rlabel metal2 8232 32200 8232 32200 0 _0283_
rlabel metal3 23576 20888 23576 20888 0 _0284_
rlabel metal2 24024 20496 24024 20496 0 _0285_
rlabel metal2 22120 20608 22120 20608 0 _0286_
rlabel metal2 14056 20048 14056 20048 0 _0287_
rlabel metal3 9912 20776 9912 20776 0 _0288_
rlabel metal3 9912 23464 9912 23464 0 _0289_
rlabel metal2 10136 31304 10136 31304 0 _0290_
rlabel metal2 17864 32872 17864 32872 0 _0291_
rlabel metal2 17640 32928 17640 32928 0 _0292_
rlabel metal3 17528 31192 17528 31192 0 _0293_
rlabel metal2 21000 34496 21000 34496 0 _0294_
rlabel metal3 24024 33488 24024 33488 0 _0295_
rlabel metal2 28280 32144 28280 32144 0 _0296_
rlabel metal2 30632 31192 30632 31192 0 _0297_
rlabel metal2 33992 29680 33992 29680 0 _0298_
rlabel metal2 32088 28616 32088 28616 0 _0299_
rlabel metal2 30408 27104 30408 27104 0 _0300_
rlabel metal2 26544 26264 26544 26264 0 _0301_
rlabel metal2 24248 20216 24248 20216 0 _0302_
rlabel metal3 20888 17864 20888 17864 0 _0303_
rlabel metal2 16408 24080 16408 24080 0 _0304_
rlabel metal3 28728 26936 28728 26936 0 _0305_
rlabel metal2 31416 32144 31416 32144 0 _0306_
rlabel metal2 35448 29904 35448 29904 0 _0307_
rlabel metal2 32536 28952 32536 28952 0 _0308_
rlabel metal2 34552 29848 34552 29848 0 _0309_
rlabel metal3 34048 28504 34048 28504 0 _0310_
rlabel metal3 35336 28616 35336 28616 0 _0311_
rlabel metal2 24696 19376 24696 19376 0 _0312_
rlabel metal2 26152 34608 26152 34608 0 _0313_
rlabel metal3 26376 23800 26376 23800 0 _0314_
rlabel metal2 31080 33376 31080 33376 0 _0315_
rlabel metal2 34216 33040 34216 33040 0 _0316_
rlabel metal2 32200 34496 32200 34496 0 _0317_
rlabel metal2 30632 33992 30632 33992 0 _0318_
rlabel metal2 18144 20104 18144 20104 0 _0319_
rlabel metal2 30688 34328 30688 34328 0 _0320_
rlabel metal2 18984 24920 18984 24920 0 _0321_
rlabel metal2 31192 36456 31192 36456 0 _0322_
rlabel metal2 23856 25592 23856 25592 0 _0323_
rlabel metal3 33096 33432 33096 33432 0 _0324_
rlabel metal2 31920 33432 31920 33432 0 _0325_
rlabel metal2 31864 35336 31864 35336 0 _0326_
rlabel metal2 32984 35616 32984 35616 0 _0327_
rlabel metal2 28056 29680 28056 29680 0 _0328_
rlabel metal2 24248 32368 24248 32368 0 _0329_
rlabel metal2 26992 32648 26992 32648 0 _0330_
rlabel metal2 27160 31696 27160 31696 0 _0331_
rlabel metal2 27608 29064 27608 29064 0 _0332_
rlabel metal2 27888 28728 27888 28728 0 _0333_
rlabel metal2 24696 29736 24696 29736 0 _0334_
rlabel metal2 27552 33432 27552 33432 0 _0335_
rlabel metal2 27608 34552 27608 34552 0 _0336_
rlabel metal2 27160 34664 27160 34664 0 _0337_
rlabel metal2 28168 36456 28168 36456 0 _0338_
rlabel metal3 23072 33208 23072 33208 0 _0339_
rlabel metal2 24584 33936 24584 33936 0 _0340_
rlabel metal2 24248 33824 24248 33824 0 _0341_
rlabel metal2 23688 33488 23688 33488 0 _0342_
rlabel metal3 24920 35000 24920 35000 0 _0343_
rlabel metal2 25704 36568 25704 36568 0 _0344_
rlabel metal2 21112 34944 21112 34944 0 _0345_
rlabel metal2 21504 34216 21504 34216 0 _0346_
rlabel metal2 21392 35896 21392 35896 0 _0347_
rlabel metal2 22008 36176 22008 36176 0 _0348_
rlabel metal2 18872 31080 18872 31080 0 _0349_
rlabel metal2 19992 31024 19992 31024 0 _0350_
rlabel metal2 20552 30464 20552 30464 0 _0351_
rlabel metal2 17080 30744 17080 30744 0 _0352_
rlabel metal2 14728 31472 14728 31472 0 _0353_
rlabel metal2 12488 30464 12488 30464 0 _0354_
rlabel metal2 15288 31304 15288 31304 0 _0355_
rlabel metal2 14392 35476 14392 35476 0 _0356_
rlabel metal3 16520 30968 16520 30968 0 _0357_
rlabel metal2 17752 30464 17752 30464 0 _0358_
rlabel metal3 19656 29512 19656 29512 0 _0359_
rlabel metal2 19432 29792 19432 29792 0 _0360_
rlabel metal2 18984 25144 18984 25144 0 _0361_
rlabel metal2 20104 29288 20104 29288 0 _0362_
rlabel metal2 17416 29008 17416 29008 0 _0363_
rlabel metal2 16968 29400 16968 29400 0 _0364_
rlabel metal3 16800 28504 16800 28504 0 _0365_
rlabel metal2 14392 27048 14392 27048 0 _0366_
rlabel metal2 14728 35896 14728 35896 0 _0367_
rlabel metal2 15176 34832 15176 34832 0 _0368_
rlabel metal2 16352 33320 16352 33320 0 _0369_
rlabel metal2 17752 34608 17752 34608 0 _0370_
rlabel metal2 18872 33432 18872 33432 0 _0371_
rlabel metal2 17080 33376 17080 33376 0 _0372_
rlabel metal2 16520 34048 16520 34048 0 _0373_
rlabel metal2 14224 36344 14224 36344 0 _0374_
rlabel metal3 16688 34888 16688 34888 0 _0375_
rlabel metal2 14728 35280 14728 35280 0 _0376_
rlabel metal2 14840 34888 14840 34888 0 _0377_
rlabel metal2 16296 35336 16296 35336 0 _0378_
rlabel metal2 18088 35056 18088 35056 0 _0379_
rlabel metal2 17752 18816 17752 18816 0 _0380_
rlabel metal2 11368 34608 11368 34608 0 _0381_
rlabel metal2 10920 33096 10920 33096 0 _0382_
rlabel metal3 10192 33544 10192 33544 0 _0383_
rlabel metal2 9240 34384 9240 34384 0 _0384_
rlabel metal2 10248 34272 10248 34272 0 _0385_
rlabel metal2 10584 35056 10584 35056 0 _0386_
rlabel metal2 12040 35728 12040 35728 0 _0387_
rlabel metal2 16744 19488 16744 19488 0 _0388_
rlabel metal2 8120 31304 8120 31304 0 _0389_
rlabel metal2 7784 32200 7784 32200 0 _0390_
rlabel metal2 8624 32648 8624 32648 0 _0391_
rlabel metal2 10696 32592 10696 32592 0 _0392_
rlabel metal2 10024 32704 10024 32704 0 _0393_
rlabel metal3 7392 33096 7392 33096 0 _0394_
rlabel metal2 6720 33320 6720 33320 0 _0395_
rlabel metal2 7000 30520 7000 30520 0 _0396_
rlabel metal3 10360 29400 10360 29400 0 _0397_
rlabel metal2 10248 29680 10248 29680 0 _0398_
rlabel metal3 6944 30072 6944 30072 0 _0399_
rlabel metal3 6160 29400 6160 29400 0 _0400_
rlabel metal2 6216 29344 6216 29344 0 _0401_
rlabel metal2 10864 27832 10864 27832 0 _0402_
rlabel metal3 10024 28056 10024 28056 0 _0403_
rlabel metal2 10472 28112 10472 28112 0 _0404_
rlabel metal2 6552 28616 6552 28616 0 _0405_
rlabel metal2 8344 22288 8344 22288 0 _0406_
rlabel metal2 8288 25480 8288 25480 0 _0407_
rlabel metal2 9464 25872 9464 25872 0 _0408_
rlabel metal2 10472 25536 10472 25536 0 _0409_
rlabel metal3 11704 25368 11704 25368 0 _0410_
rlabel metal2 9576 20384 9576 20384 0 _0411_
rlabel metal2 10136 24976 10136 24976 0 _0412_
rlabel metal2 11592 25816 11592 25816 0 _0413_
rlabel metal2 12152 26208 12152 26208 0 _0414_
rlabel metal2 13608 26264 13608 26264 0 _0415_
rlabel metal2 8064 24808 8064 24808 0 _0416_
rlabel metal2 7336 26096 7336 26096 0 _0417_
rlabel metal2 5656 25816 5656 25816 0 _0418_
rlabel metal2 6328 25480 6328 25480 0 _0419_
rlabel metal2 8904 20552 8904 20552 0 _0420_
rlabel metal3 8064 19432 8064 19432 0 _0421_
rlabel metal2 8904 19712 8904 19712 0 _0422_
rlabel metal3 7784 22456 7784 22456 0 _0423_
rlabel metal2 7112 21168 7112 21168 0 _0424_
rlabel metal3 8176 19992 8176 19992 0 _0425_
rlabel metal2 4536 19264 4536 19264 0 _0426_
rlabel metal2 5376 19208 5376 19208 0 _0427_
rlabel metal2 8008 21224 8008 21224 0 _0428_
rlabel metal2 8568 22288 8568 22288 0 _0429_
rlabel metal2 8792 21896 8792 21896 0 _0430_
rlabel metal2 4536 20888 4536 20888 0 _0431_
rlabel metal2 5320 20776 5320 20776 0 _0432_
rlabel metal2 9296 18424 9296 18424 0 _0433_
rlabel metal2 12488 16464 12488 16464 0 _0434_
rlabel metal3 13216 19208 13216 19208 0 _0435_
rlabel metal2 13496 17920 13496 17920 0 _0436_
rlabel metal2 11144 17472 11144 17472 0 _0437_
rlabel metal2 10360 17304 10360 17304 0 _0438_
rlabel metal2 8904 17976 8904 17976 0 _0439_
rlabel metal2 9688 17640 9688 17640 0 _0440_
rlabel metal2 14056 18928 14056 18928 0 _0441_
rlabel metal2 13608 18368 13608 18368 0 _0442_
rlabel metal2 13160 19040 13160 19040 0 _0443_
rlabel metal2 14280 17808 14280 17808 0 _0444_
rlabel metal2 11816 17024 11816 17024 0 _0445_
rlabel metal3 13216 16856 13216 16856 0 _0446_
rlabel metal2 17752 21056 17752 21056 0 _0447_
rlabel metal2 17416 20328 17416 20328 0 _0448_
rlabel metal3 18592 22120 18592 22120 0 _0449_
rlabel metal2 18088 22624 18088 22624 0 _0450_
rlabel metal2 15736 20832 15736 20832 0 _0451_
rlabel metal2 17864 20272 17864 20272 0 _0452_
rlabel metal2 17024 19208 17024 19208 0 _0453_
rlabel metal3 17192 18424 17192 18424 0 _0454_
rlabel metal2 14728 21952 14728 21952 0 _0455_
rlabel metal2 17640 22064 17640 22064 0 _0456_
rlabel metal3 16912 22232 16912 22232 0 _0457_
rlabel metal2 17416 22792 17416 22792 0 _0458_
rlabel metal2 17752 24108 17752 24108 0 _0459_
rlabel metal3 24080 20552 24080 20552 0 _0460_
rlabel metal2 22232 23520 22232 23520 0 _0461_
rlabel metal2 22736 24808 22736 24808 0 _0462_
rlabel metal2 21056 24696 21056 24696 0 _0463_
rlabel metal2 21056 24920 21056 24920 0 _0464_
rlabel metal2 21560 25928 21560 25928 0 _0465_
rlabel metal2 22456 26320 22456 26320 0 _0466_
rlabel metal2 22960 28056 22960 28056 0 _0467_
rlabel metal2 23576 27888 23576 27888 0 _0468_
rlabel metal2 20664 21672 20664 21672 0 _0469_
rlabel metal2 21728 22456 21728 22456 0 _0470_
rlabel metal2 21224 23408 21224 23408 0 _0471_
rlabel metal2 21000 23464 21000 23464 0 _0472_
rlabel metal2 21784 24360 21784 24360 0 _0473_
rlabel metal2 19432 24752 19432 24752 0 _0474_
rlabel metal3 25536 23128 25536 23128 0 _0475_
rlabel metal2 26096 19208 26096 19208 0 _0476_
rlabel metal3 25760 19992 25760 19992 0 _0477_
rlabel metal2 26600 19432 26600 19432 0 _0478_
rlabel metal3 25592 19096 25592 19096 0 _0479_
rlabel metal2 23800 20048 23800 20048 0 _0480_
rlabel metal2 29064 22624 29064 22624 0 _0481_
rlabel metal2 27384 23520 27384 23520 0 _0482_
rlabel metal2 27888 21672 27888 21672 0 _0483_
rlabel metal2 27160 24360 27160 24360 0 _0484_
rlabel metal2 26152 24752 26152 24752 0 _0485_
rlabel metal2 34664 24360 34664 24360 0 _0486_
rlabel metal2 35952 24920 35952 24920 0 _0487_
rlabel metal2 32200 24976 32200 24976 0 _0488_
rlabel metal2 31528 24864 31528 24864 0 _0489_
rlabel metal2 30968 20944 30968 20944 0 _0490_
rlabel metal3 29960 21000 29960 21000 0 _0491_
rlabel metal3 30520 21784 30520 21784 0 _0492_
rlabel metal2 29736 25760 29736 25760 0 _0493_
rlabel metal2 33992 24472 33992 24472 0 _0494_
rlabel metal2 31192 20048 31192 20048 0 _0495_
rlabel metal2 31528 21392 31528 21392 0 _0496_
rlabel metal2 32536 26432 32536 26432 0 _0497_
rlabel metal2 33208 18928 33208 18928 0 _0498_
rlabel metal3 33992 20776 33992 20776 0 _0499_
rlabel metal2 33096 21056 33096 21056 0 _0500_
rlabel metal2 33432 20216 33432 20216 0 _0501_
rlabel metal2 34776 19488 34776 19488 0 _0502_
rlabel metal3 33264 21560 33264 21560 0 _0503_
rlabel metal2 32816 21336 32816 21336 0 _0504_
rlabel metal3 33544 21784 33544 21784 0 _0505_
rlabel metal2 25480 10584 25480 10584 0 _0506_
rlabel metal3 21980 13048 21980 13048 0 _0507_
rlabel metal2 25256 10920 25256 10920 0 _0508_
rlabel metal2 25928 10416 25928 10416 0 _0509_
rlabel metal3 21224 14504 21224 14504 0 _0510_
rlabel metal3 26600 13552 26600 13552 0 _0511_
rlabel metal2 28504 8400 28504 8400 0 _0512_
rlabel metal3 32704 9128 32704 9128 0 _0513_
rlabel metal2 33040 15512 33040 15512 0 _0514_
rlabel metal2 35672 12880 35672 12880 0 _0515_
rlabel metal2 33992 15288 33992 15288 0 _0516_
rlabel metal3 35280 15064 35280 15064 0 _0517_
rlabel metal2 33992 9744 33992 9744 0 _0518_
rlabel metal3 31864 9016 31864 9016 0 _0519_
rlabel metal2 30296 8960 30296 8960 0 _0520_
rlabel metal2 28616 8064 28616 8064 0 _0521_
rlabel metal2 28280 8400 28280 8400 0 _0522_
rlabel metal2 27776 9128 27776 9128 0 _0523_
rlabel metal2 27384 9912 27384 9912 0 _0524_
rlabel metal2 33096 12544 33096 12544 0 _0525_
rlabel metal2 27944 12488 27944 12488 0 _0526_
rlabel metal3 33152 13160 33152 13160 0 _0527_
rlabel metal2 34104 12152 34104 12152 0 _0528_
rlabel metal2 23240 9464 23240 9464 0 _0529_
rlabel metal2 32648 15736 32648 15736 0 _0530_
rlabel metal2 30744 12600 30744 12600 0 _0531_
rlabel metal2 31080 11984 31080 11984 0 _0532_
rlabel metal2 30408 11088 30408 11088 0 _0533_
rlabel metal2 27832 11368 27832 11368 0 _0534_
rlabel metal3 28448 12936 28448 12936 0 _0535_
rlabel metal2 26600 14168 26600 14168 0 _0536_
rlabel metal2 28504 13216 28504 13216 0 _0537_
rlabel metal3 28896 13160 28896 13160 0 _0538_
rlabel metal2 26488 13160 26488 13160 0 _0539_
rlabel metal2 26376 13608 26376 13608 0 _0540_
rlabel metal2 27048 11144 27048 11144 0 _0541_
rlabel metal2 24808 9856 24808 9856 0 _0542_
rlabel metal2 22904 12992 22904 12992 0 _0543_
rlabel metal2 25144 10640 25144 10640 0 _0544_
rlabel metal2 26824 9408 26824 9408 0 _0545_
rlabel metal3 29680 9240 29680 9240 0 _0546_
rlabel metal2 28840 11368 28840 11368 0 _0547_
rlabel metal2 30408 9912 30408 9912 0 _0548_
rlabel metal3 30464 9576 30464 9576 0 _0549_
rlabel metal2 33768 9296 33768 9296 0 _0550_
rlabel metal3 31304 11200 31304 11200 0 _0551_
rlabel metal3 31136 10808 31136 10808 0 _0552_
rlabel metal2 30520 11480 30520 11480 0 _0553_
rlabel metal2 33096 8960 33096 8960 0 _0554_
rlabel metal2 33432 9464 33432 9464 0 _0555_
rlabel metal3 33376 10024 33376 10024 0 _0556_
rlabel metal2 33096 11032 33096 11032 0 _0557_
rlabel metal2 32480 13160 32480 13160 0 _0558_
rlabel metal2 33264 12936 33264 12936 0 _0559_
rlabel metal2 33432 13328 33432 13328 0 _0560_
rlabel metal2 32760 11592 32760 11592 0 _0561_
rlabel metal3 34552 11256 34552 11256 0 _0562_
rlabel metal2 35784 11368 35784 11368 0 _0563_
rlabel metal2 30296 14056 30296 14056 0 _0564_
rlabel metal2 30184 12936 30184 12936 0 _0565_
rlabel metal2 29848 13048 29848 13048 0 _0566_
rlabel metal2 29288 13160 29288 13160 0 _0567_
rlabel metal2 34104 13216 34104 13216 0 _0568_
rlabel metal3 35392 12936 35392 12936 0 _0569_
rlabel metal2 21112 13216 21112 13216 0 _0570_
rlabel metal2 21112 14000 21112 14000 0 _0571_
rlabel metal2 19600 8120 19600 8120 0 _0572_
rlabel metal2 19600 11256 19600 11256 0 _0573_
rlabel metal2 17528 11312 17528 11312 0 _0574_
rlabel metal2 26824 14112 26824 14112 0 _0575_
rlabel metal3 26040 13272 26040 13272 0 _0576_
rlabel metal2 31976 15792 31976 15792 0 _0577_
rlabel metal3 33936 15960 33936 15960 0 _0578_
rlabel metal3 31192 15176 31192 15176 0 _0579_
rlabel metal2 27440 13608 27440 13608 0 _0580_
rlabel metal2 27832 14672 27832 14672 0 _0581_
rlabel metal2 14728 9520 14728 9520 0 _0582_
rlabel metal2 25480 17248 25480 17248 0 _0583_
rlabel metal3 16072 15176 16072 15176 0 _0584_
rlabel metal3 38920 10696 38920 10696 0 _0585_
rlabel metal2 21448 18928 21448 18928 0 _0586_
rlabel metal2 20776 25032 20776 25032 0 _0587_
rlabel metal2 25928 18256 25928 18256 0 _0588_
rlabel metal2 11256 11424 11256 11424 0 _0589_
rlabel metal2 11368 12320 11368 12320 0 _0590_
rlabel metal2 13160 10976 13160 10976 0 _0591_
rlabel metal3 10136 10024 10136 10024 0 _0592_
rlabel metal2 5656 13384 5656 13384 0 _0593_
rlabel metal3 8008 14392 8008 14392 0 _0594_
rlabel metal2 22344 19152 22344 19152 0 clknet_0_clock
rlabel metal2 2296 14896 2296 14896 0 clknet_2_0__leaf_clock
rlabel metal2 16632 25536 16632 25536 0 clknet_2_1__leaf_clock
rlabel metal3 20944 16072 20944 16072 0 clknet_2_2__leaf_clock
rlabel metal2 19544 37408 19544 37408 0 clknet_2_3__leaf_clock
rlabel metal2 18592 20216 18592 20216 0 clock
rlabel metal2 16856 854 16856 854 0 logisim_clock_tree_0_out
rlabel metal2 7616 13160 7616 13160 0 manchester_baby_instance.BASE_0.s_countReg\[0\]
rlabel metal2 7336 13720 7336 13720 0 manchester_baby_instance.BASE_0.s_countReg\[1\]
rlabel metal2 7224 13720 7224 13720 0 manchester_baby_instance.BASE_0.s_countReg\[2\]
rlabel metal3 8232 12824 8232 12824 0 manchester_baby_instance.BASE_0.s_tickNext
rlabel metal3 11480 13048 11480 13048 0 manchester_baby_instance.BASE_0.s_tickReg
rlabel metal2 14392 11256 14392 11256 0 manchester_baby_instance.BASE_1.s_bufferRegs\[0\]
rlabel metal2 11424 9912 11424 9912 0 manchester_baby_instance.BASE_1.s_counterValue
rlabel metal2 13944 10640 13944 10640 0 manchester_baby_instance.BASE_1.s_derivedClock
rlabel metal2 34440 15204 34440 15204 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\]
rlabel metal2 38360 10976 38360 10976 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\]
rlabel metal2 30632 12096 30632 12096 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\]
rlabel metal2 28280 13552 28280 13552 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\]
rlabel metal2 27048 8008 27048 8008 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\]
rlabel metal2 20384 17640 20384 17640 0 manchester_baby_instance.CIRCUIT_0.Acc.tick
rlabel metal2 18200 8232 18200 8232 0 manchester_baby_instance.CIRCUIT_0.GATES_13.result
rlabel metal2 33208 17248 33208 17248 0 manchester_baby_instance.CIRCUIT_0.IR.q\[0\]
rlabel metal2 25480 15288 25480 15288 0 manchester_baby_instance.CIRCUIT_0.IR.q\[13\]
rlabel metal3 19768 16072 19768 16072 0 manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
rlabel metal3 17864 16296 17864 16296 0 manchester_baby_instance.CIRCUIT_0.IR.q\[15\]
rlabel metal2 34160 15960 34160 15960 0 manchester_baby_instance.CIRCUIT_0.IR.q\[1\]
rlabel metal2 30296 15792 30296 15792 0 manchester_baby_instance.CIRCUIT_0.IR.q\[2\]
rlabel metal2 25704 9856 25704 9856 0 manchester_baby_instance.CIRCUIT_0.IR.q\[3\]
rlabel metal2 27160 16688 27160 16688 0 manchester_baby_instance.CIRCUIT_0.IR.q\[4\]
rlabel metal2 20776 10920 20776 10920 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
rlabel metal2 22232 12936 22232 12936 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
rlabel metal2 22904 10192 22904 10192 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\]
rlabel metal2 22008 13104 22008 13104 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[0\]
rlabel metal2 18872 7728 18872 7728 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[1\]
rlabel metal2 18760 10864 18760 10864 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[2\]
rlabel metal2 39256 15176 39256 15176 0 net1
rlabel metal3 9632 34664 9632 34664 0 net10
rlabel metal2 11928 34496 11928 34496 0 net11
rlabel metal2 39704 12600 39704 12600 0 net12
rlabel metal2 15960 35952 15960 35952 0 net13
rlabel metal2 15456 35112 15456 35112 0 net14
rlabel metal2 18648 35560 18648 35560 0 net15
rlabel metal3 19544 31640 19544 31640 0 net16
rlabel metal2 23016 35056 23016 35056 0 net17
rlabel metal2 23576 35896 23576 35896 0 net18
rlabel metal3 26824 33824 26824 33824 0 net19
rlabel metal2 2296 17976 2296 17976 0 net2
rlabel metal2 28056 32760 28056 32760 0 net20
rlabel metal2 35000 31640 35000 31640 0 net21
rlabel metal2 39256 30912 39256 30912 0 net22
rlabel metal3 39928 19264 39928 19264 0 net23
rlabel metal2 39928 31472 39928 31472 0 net24
rlabel metal2 39928 28840 39928 28840 0 net25
rlabel metal3 28504 19096 28504 19096 0 net26
rlabel metal2 26824 17640 26824 17640 0 net27
rlabel metal2 39256 21672 39256 21672 0 net28
rlabel metal2 26712 20944 26712 20944 0 net29
rlabel metal2 11032 19152 11032 19152 0 net3
rlabel metal2 39928 22680 39928 22680 0 net30
rlabel metal2 2296 20384 2296 20384 0 net31
rlabel metal2 3192 20216 3192 20216 0 net32
rlabel metal2 23352 18424 23352 18424 0 net33
rlabel metal2 17752 8120 17752 8120 0 net34
rlabel metal2 39144 16576 39144 16576 0 net35
rlabel metal2 39032 16576 39032 16576 0 net36
rlabel metal2 31640 15792 31640 15792 0 net37
rlabel metal2 25368 14448 25368 14448 0 net38
rlabel metal2 39032 15008 39032 15008 0 net39
rlabel metal2 6216 21616 6216 21616 0 net4
rlabel metal2 39144 21952 39144 21952 0 net40
rlabel metal2 2968 16128 2968 16128 0 net41
rlabel metal2 10024 17248 10024 17248 0 net42
rlabel metal2 2856 22232 2856 22232 0 net43
rlabel metal2 5768 19152 5768 19152 0 net44
rlabel metal2 2856 25592 2856 25592 0 net45
rlabel metal2 2968 25536 2968 25536 0 net46
rlabel metal2 2968 28672 2968 28672 0 net47
rlabel metal2 2856 30464 2856 30464 0 net48
rlabel metal2 8680 36400 8680 36400 0 net49
rlabel metal2 3192 18368 3192 18368 0 net5
rlabel metal2 12600 36736 12600 36736 0 net50
rlabel metal2 34160 19992 34160 19992 0 net51
rlabel metal2 17696 35672 17696 35672 0 net52
rlabel via2 16184 36904 16184 36904 0 net53
rlabel metal3 17416 28728 17416 28728 0 net54
rlabel metal2 21784 30184 21784 30184 0 net55
rlabel metal2 23240 37744 23240 37744 0 net56
rlabel metal2 25368 37184 25368 37184 0 net57
rlabel metal2 29736 37464 29736 37464 0 net58
rlabel metal2 26768 30968 26768 30968 0 net59
rlabel metal2 2072 24976 2072 24976 0 net6
rlabel metal3 36064 36680 36064 36680 0 net60
rlabel metal2 32760 37016 32760 37016 0 net61
rlabel metal2 36568 25984 36568 25984 0 net62
rlabel via2 37464 28728 37464 28728 0 net63
rlabel metal2 38696 13384 38696 13384 0 net64
rlabel metal2 31472 24584 31472 24584 0 net65
rlabel metal3 38836 23912 38836 23912 0 net66
rlabel metal2 39032 21000 39032 21000 0 net67
rlabel metal3 19600 25704 19600 25704 0 net68
rlabel metal2 23800 24696 23800 24696 0 net69
rlabel metal3 2296 23856 2296 23856 0 net7
rlabel metal2 2856 23240 2856 23240 0 net70
rlabel metal2 2744 19264 2744 19264 0 net71
rlabel metal3 21448 3416 21448 3416 0 net72
rlabel metal2 18592 11144 18592 11144 0 net73
rlabel metal2 14728 12656 14728 12656 0 net74
rlabel metal2 2072 29176 2072 29176 0 net8
rlabel metal2 7784 31696 7784 31696 0 net9
rlabel metal2 40040 17304 40040 17304 0 ram_addr_o[0]
rlabel metal2 39816 16520 39816 16520 0 ram_addr_o[1]
rlabel metal2 40152 15736 40152 15736 0 ram_addr_o[2]
rlabel metal2 26264 854 26264 854 0 ram_addr_o[3]
rlabel metal2 39816 15008 39816 15008 0 ram_addr_o[4]
rlabel metal2 40264 14336 40264 14336 0 ram_data_i[0]
rlabel metal3 1246 17528 1246 17528 0 ram_data_i[10]
rlabel metal3 2072 18144 2072 18144 0 ram_data_i[11]
rlabel metal3 1358 22232 1358 22232 0 ram_data_i[12]
rlabel metal2 2632 17136 2632 17136 0 ram_data_i[13]
rlabel metal2 1736 24472 1736 24472 0 ram_data_i[14]
rlabel metal2 1736 23632 1736 23632 0 ram_data_i[15]
rlabel metal2 1736 29176 1736 29176 0 ram_data_i[16]
rlabel metal2 1736 31248 1736 31248 0 ram_data_i[17]
rlabel metal2 9464 39942 9464 39942 0 ram_data_i[18]
rlabel metal2 11480 39942 11480 39942 0 ram_data_i[19]
rlabel metal3 40754 12824 40754 12824 0 ram_data_i[1]
rlabel metal2 16744 37800 16744 37800 0 ram_data_i[20]
rlabel metal2 16856 39942 16856 39942 0 ram_data_i[21]
rlabel metal2 18200 39942 18200 39942 0 ram_data_i[22]
rlabel metal2 18872 39942 18872 39942 0 ram_data_i[23]
rlabel metal2 24024 37520 24024 37520 0 ram_data_i[24]
rlabel metal2 23576 39942 23576 39942 0 ram_data_i[25]
rlabel metal2 27384 35840 27384 35840 0 ram_data_i[26]
rlabel metal2 30296 37352 30296 37352 0 ram_data_i[27]
rlabel metal2 31640 39942 31640 39942 0 ram_data_i[28]
rlabel metal3 40418 31640 40418 31640 0 ram_data_i[29]
rlabel metal2 40264 20440 40264 20440 0 ram_data_i[2]
rlabel metal3 40754 30968 40754 30968 0 ram_data_i[30]
rlabel metal2 40264 28448 40264 28448 0 ram_data_i[31]
rlabel metal2 40264 18984 40264 18984 0 ram_data_i[3]
rlabel metal2 25816 2520 25816 2520 0 ram_data_i[4]
rlabel metal2 39592 22344 39592 22344 0 ram_data_i[5]
rlabel metal2 21560 39942 21560 39942 0 ram_data_i[6]
rlabel metal2 40264 23016 40264 23016 0 ram_data_i[7]
rlabel metal2 1736 20832 1736 20832 0 ram_data_i[8]
rlabel metal2 2632 20384 2632 20384 0 ram_data_i[9]
rlabel metal2 40040 22344 40040 22344 0 ram_data_o[0]
rlabel metal3 1414 15512 1414 15512 0 ram_data_o[10]
rlabel metal3 1470 16184 1470 16184 0 ram_data_o[11]
rlabel metal3 1470 21560 1470 21560 0 ram_data_o[12]
rlabel metal3 1414 18872 1414 18872 0 ram_data_o[13]
rlabel metal3 1358 25592 1358 25592 0 ram_data_o[14]
rlabel metal3 1470 24920 1470 24920 0 ram_data_o[15]
rlabel metal3 1470 28280 1470 28280 0 ram_data_o[16]
rlabel metal3 1470 30296 1470 30296 0 ram_data_o[17]
rlabel metal2 9800 38360 9800 38360 0 ram_data_o[18]
rlabel metal2 13160 38416 13160 38416 0 ram_data_o[19]
rlabel metal2 40040 19712 40040 19712 0 ram_data_o[1]
rlabel metal3 18872 38248 18872 38248 0 ram_data_o[20]
rlabel metal2 14840 39746 14840 39746 0 ram_data_o[21]
rlabel metal3 16800 37464 16800 37464 0 ram_data_o[22]
rlabel metal2 21112 39592 21112 39592 0 ram_data_o[23]
rlabel metal2 22904 39690 22904 39690 0 ram_data_o[24]
rlabel metal2 26376 38360 26376 38360 0 ram_data_o[25]
rlabel metal2 30408 38192 30408 38192 0 ram_data_o[26]
rlabel metal2 26264 39914 26264 39914 0 ram_data_o[27]
rlabel metal2 34384 38136 34384 38136 0 ram_data_o[28]
rlabel metal2 32536 39480 32536 39480 0 ram_data_o[29]
rlabel metal2 40152 25872 40152 25872 0 ram_data_o[2]
rlabel metal2 40152 29120 40152 29120 0 ram_data_o[30]
rlabel metal2 40040 13552 40040 13552 0 ram_data_o[31]
rlabel metal2 39816 25088 39816 25088 0 ram_data_o[3]
rlabel metal2 40040 23800 40040 23800 0 ram_data_o[4]
rlabel metal2 40152 21168 40152 21168 0 ram_data_o[5]
rlabel metal2 20216 39746 20216 39746 0 ram_data_o[6]
rlabel metal2 24528 39592 24528 39592 0 ram_data_o[7]
rlabel metal3 1358 22904 1358 22904 0 ram_data_o[8]
rlabel metal3 1358 19544 1358 19544 0 ram_data_o[9]
rlabel metal2 21896 3640 21896 3640 0 ram_rw_en_o
rlabel metal2 22904 2058 22904 2058 0 reset_i
rlabel metal3 18536 3640 18536 3640 0 stop_lamp_o
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
