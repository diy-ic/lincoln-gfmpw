module manchester_baby (clock,
    logisim_clock_tree_0_out,
    ram_rw_en_o,
    reset_i,
    stop_lamp_o,
    vdd,
    vss,
    ram_addr_o,
    ram_data_i,
    ram_data_o);
 input clock;
 output logisim_clock_tree_0_out;
 output ram_rw_en_o;
 input reset_i;
 output stop_lamp_o;
 input vdd;
 input vss;
 output [4:0] ram_addr_o;
 input [31:0] ram_data_i;
 output [31:0] ram_data_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire clknet_0_clock;
 wire clknet_2_0__leaf_clock;
 wire clknet_2_1__leaf_clock;
 wire clknet_2_2__leaf_clock;
 wire clknet_2_3__leaf_clock;
 wire \manchester_baby_instance.BASE_0.s_countReg[0] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[1] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[2] ;
 wire \manchester_baby_instance.BASE_0.s_tickNext ;
 wire \manchester_baby_instance.BASE_0.s_tickReg ;
 wire \manchester_baby_instance.BASE_1.s_bufferRegs[0] ;
 wire \manchester_baby_instance.BASE_1.s_counterValue ;
 wire \manchester_baby_instance.BASE_1.s_derivedClock ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ;
 wire \manchester_baby_instance.CIRCUIT_0.Acc.tick ;
 wire \manchester_baby_instance.CIRCUIT_0.GATES_13.result ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[13] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[14] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[15] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[2] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[3] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[4] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[2] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net8;
 wire net9;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0605__I (.I(_0108_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0606__A2 (.I(_0109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0607__A2 (.I(_0109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0609__A2 (.I(_0109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0610__A2 (.I(_0109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0612__A1 (.I(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0612__A2 (.I(_0108_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0613__A2 (.I(_0109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0614__I (.I(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0615__A2 (.I(_0109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0616__A2 (.I(_0109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0618__I0 (.I(_0117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0618__S (.I(_0108_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0621__I0 (.I(_0119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0621__S (.I(_0108_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0623__I (.I(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0624__A2 (.I(_0109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0625__A2 (.I(_0109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0627__A2 (.I(_0108_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0628__A2 (.I(_0109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0670__A1 (.I(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0677__I (.I(net71),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0678__I (.I(net31),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0680__A1 (.I(net70),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0680__B2 (.I(net71),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0687__I (.I(net30),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0689__I (.I(net29),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0694__A1 (.I(_0117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0696__A1 (.I(_0117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0696__C (.I(_0119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0698__A1 (.I(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0700__A1 (.I(_0119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0701__A1 (.I(_0117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0704__A1 (.I(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0719__A1 (.I(net70),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0726__A1 (.I(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0729__A1 (.I(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0780__A1 (.I(net64),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0788__A1 (.I(_0117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0788__A3 (.I(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0789__A1 (.I(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0790__A1 (.I(net29),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0790__A2 (.I(net30),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0791__A1 (.I(net31),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0792__A1 (.I(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0804__A1 (.I(_0126_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0804__B1 (.I(_0281_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0807__A1 (.I(_0301_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0807__A2 (.I(_0302_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0809__I1 (.I(net64),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0809__S (.I(_0304_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0813__A1 (.I(_0301_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0815__A1 (.I(_0281_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0816__S (.I(_0304_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0819__I (.I(_0312_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0820__I (.I(_0302_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0825__I (.I(_0301_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0826__A1 (.I(_0314_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0826__B2 (.I(_0319_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0827__I (.I(_0312_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0828__A2 (.I(_0321_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0829__A1 (.I(_0313_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0830__I (.I(_0301_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0833__A1 (.I(_0323_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0833__B2 (.I(_0314_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0834__A2 (.I(_0321_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0835__A1 (.I(_0313_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0841__A1 (.I(_0281_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0841__B2 (.I(_0126_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0842__S (.I(_0304_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0846__A1 (.I(_0323_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0846__B2 (.I(_0314_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0847__A2 (.I(_0321_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0848__A1 (.I(_0313_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0853__A1 (.I(_0314_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0853__B2 (.I(_0319_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0854__A2 (.I(_0321_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0855__A1 (.I(_0313_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0858__A1 (.I(_0314_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0858__B2 (.I(_0319_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0859__A2 (.I(_0321_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0860__A1 (.I(_0313_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0872__A1 (.I(_0314_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0872__B2 (.I(_0319_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0874__A2 (.I(_0361_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0875__A1 (.I(_0313_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0878__A1 (.I(_0281_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0878__B2 (.I(_0126_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0879__S (.I(_0312_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0886__A1 (.I(_0302_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0887__A1 (.I(_0126_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0888__S (.I(_0312_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0892__A1 (.I(_0126_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0893__A1 (.I(_0314_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0894__A2 (.I(_0361_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0895__A1 (.I(_0313_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0896__I (.I(_0302_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0902__A1 (.I(_0380_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0902__B2 (.I(_0319_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0903__A2 (.I(_0361_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0904__A1 (.I(_0313_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0905__I (.I(_0312_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0909__A1 (.I(_0301_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0911__A1 (.I(_0314_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0912__A2 (.I(_0361_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0913__A1 (.I(_0388_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0918__A1 (.I(_0380_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0918__B2 (.I(_0319_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0919__A2 (.I(_0361_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0920__A1 (.I(_0388_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0923__A1 (.I(_0323_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0923__B2 (.I(_0314_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0924__A2 (.I(_0361_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0925__A1 (.I(_0388_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0933__A1 (.I(_0281_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0934__A1 (.I(_0323_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0935__A2 (.I(_0361_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0936__A1 (.I(_0388_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0939__A1 (.I(_0380_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0939__B2 (.I(_0319_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0940__A2 (.I(_0361_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0941__A1 (.I(_0388_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0943__B (.I(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0948__A1 (.I(_0380_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0948__B2 (.I(_0319_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0949__A2 (.I(_0361_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0950__A1 (.I(_0388_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0953__A1 (.I(_0126_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0954__A1 (.I(_0380_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0955__A2 (.I(_0361_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0956__A1 (.I(_0388_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0963__A1 (.I(_0380_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0963__B2 (.I(_0319_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0964__A2 (.I(_0304_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0965__A1 (.I(_0388_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0966__A1 (.I(net31),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0967__A1 (.I(_0281_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0969__A1 (.I(_0126_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0971__A2 (.I(_0304_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0972__A1 (.I(_0388_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0973__A1 (.I(net31),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0975__A1 (.I(net70),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0979__A1 (.I(_0380_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0979__B2 (.I(_0319_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0980__A1 (.I(net71),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0980__A2 (.I(_0304_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0981__A1 (.I(_0388_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0982__A1 (.I(net31),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0983__A1 (.I(_0281_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0985__B2 (.I(_0323_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0986__A1 (.I(net70),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0986__A2 (.I(_0304_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0987__A1 (.I(_0321_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0989__A1 (.I(net29),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0995__A1 (.I(_0380_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0995__B2 (.I(_0323_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0996__A2 (.I(_0304_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0997__A1 (.I(_0321_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0998__A1 (.I(net29),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0999__A1 (.I(_0281_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1001__A1 (.I(_0301_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1003__A2 (.I(_0304_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1004__A1 (.I(_0321_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1007__A1 (.I(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1008__A1 (.I(_0302_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1009__A1 (.I(_0126_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1010__S (.I(_0312_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1013__A1 (.I(_0301_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1014__A1 (.I(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1015__B2 (.I(_0314_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1016__A2 (.I(_0304_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1017__A1 (.I(_0321_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1020__A1 (.I(_0119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1022__A1 (.I(_0119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1022__A2 (.I(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1023__A1 (.I(_0302_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1024__A1 (.I(_0117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1025__A1 (.I(_0323_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1025__C (.I(_0312_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1026__A2 (.I(_0313_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1028__A1 (.I(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1028__B (.I(_0119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1030__A1 (.I(_0323_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1030__B2 (.I(_0380_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1030__C (.I(_0312_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1031__A2 (.I(_0313_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1034__A1 (.I(_0323_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1035__A1 (.I(_0281_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1036__S (.I(_0312_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1039__A2 (.I(_0380_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1040__A2 (.I(_0323_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1040__B (.I(_0312_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1041__A2 (.I(_0321_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1048__A1 (.I(_0117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1049__A1 (.I(_0119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1051__A1 (.I(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1052__A1 (.I(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1055__A1 (.I(_0119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1057__A1 (.I(_0117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1059__A1 (.I(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1063__A1 (.I(net64),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1073__A1 (.I(net64),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1077__A1 (.I(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1083__A1 (.I(_0117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1085__A1 (.I(_0117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1088__A1 (.I(_0119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1090__A1 (.I(_0119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1097__A1 (.I(net64),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1101__A1 (.I(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1104__A1 (.I(net64),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1137__I (.I(_0584_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1138__I (.I(_0585_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1139__I (.I(_0585_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1140__I (.I(_0585_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1141__I (.I(_0585_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1142__I (.I(_0585_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1143__I (.I(_0585_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1144__I (.I(_0585_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1145__I (.I(_0585_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1146__I (.I(_0585_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1147__I (.I(_0585_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1149__I (.I(_0586_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1150__I (.I(_0586_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1151__I (.I(_0586_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1152__I (.I(_0586_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1153__I (.I(_0586_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1154__I (.I(_0586_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1155__I (.I(_0586_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1156__I (.I(_0586_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1157__I (.I(_0586_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1158__I (.I(_0586_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1160__I (.I(_0587_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1161__I (.I(_0587_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1162__I (.I(_0587_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1163__I (.I(_0587_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1164__I (.I(_0587_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1165__I (.I(_0587_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1166__I (.I(_0587_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1167__I (.I(_0587_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1168__I (.I(_0587_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1169__I (.I(_0587_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1171__I (.I(_0588_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1172__I (.I(_0588_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1173__I (.I(_0588_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1174__I (.I(_0588_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1175__I (.I(_0588_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1176__I (.I(_0588_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1177__I (.I(_0588_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1178__I (.I(_0588_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1179__I (.I(_0588_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1180__I (.I(_0588_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1181__I (.I(_0584_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1182__I (.I(_0584_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1183__I (.I(_0584_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1184__I (.I(_0584_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1185__I (.I(_0584_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1190__I (.I(_0584_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1191__I (.I(_0584_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1192__I (.I(_0584_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1193__I (.I(_0584_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1201__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1202__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1203__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1204__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1205__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1206__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1207__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1208__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1209__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1210__CLK (.I(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1211__CLK (.I(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1212__CLK (.I(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1213__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1214__CLK (.I(clknet_2_1__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1215__CLK (.I(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1216__CLK (.I(clknet_2_1__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1217__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1218__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1219__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1220__CLK (.I(clknet_2_1__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1221__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1222__CLK (.I(clknet_2_1__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1223__CLK (.I(clknet_2_1__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1224__CLK (.I(clknet_2_1__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1225__CLK (.I(clknet_2_1__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1226__CLK (.I(clknet_2_1__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1227__CLK (.I(clknet_2_1__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1228__CLK (.I(clknet_2_1__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1229__CLK (.I(clknet_2_1__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1230__CLK (.I(clknet_2_1__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1231__CLK (.I(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1232__CLK (.I(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1233__CLK (.I(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1234__CLK (.I(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1235__CLK (.I(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1236__CLK (.I(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1237__CLK (.I(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1238__CLK (.I(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1239__CLK (.I(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1240__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1241__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1242__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1243__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1244__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1245__CLK (.I(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1246__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1247__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1248__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1252__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1253__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1254__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1255__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1256__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1257__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1258__CLK (.I(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clock_I (.I(clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_clock_I (.I(clknet_0_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_clock_I (.I(clknet_0_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_clock_I (.I(clknet_0_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_clock_I (.I(clknet_0_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(ram_data_i[18]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(ram_data_i[19]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(ram_data_i[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(ram_data_i[20]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(ram_data_i[21]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(ram_data_i[22]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(ram_data_i[23]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(ram_data_i[24]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(ram_data_i[25]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(ram_data_i[26]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(ram_data_i[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(ram_data_i[27]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(ram_data_i[28]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(ram_data_i[29]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(ram_data_i[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(ram_data_i[30]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(ram_data_i[31]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(ram_data_i[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(ram_data_i[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(ram_data_i[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(ram_data_i[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(ram_data_i[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(ram_data_i[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(ram_data_i[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(ram_data_i[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(reset_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(ram_data_i[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(ram_data_i[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(ram_data_i[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(ram_data_i[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(ram_data_i[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(ram_data_i[16]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(ram_data_i[17]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output64_I (.I(net64),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output70_I (.I(net70),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output71_I (.I(net71),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_180 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_175 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_175 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0595_ (.A1(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .A2(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .ZN(_0101_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0596_ (.A1(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .A2(_0101_),
    .ZN(_0102_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0597_ (.A1(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .A2(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .ZN(_0103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0598_ (.A1(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .A2(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .ZN(_0104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0599_ (.I(net73),
    .ZN(_0105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0600_ (.A1(_0102_),
    .A2(_0103_),
    .A3(_0104_),
    .B(_0105_),
    .ZN(_0096_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0601_ (.I(net7),
    .ZN(_0106_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _0602_ (.I(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .ZN(_0107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _0603_ (.I(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .ZN(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0604_ (.A1(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .A2(_0107_),
    .A3(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .A4(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ),
    .ZN(_0108_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0605_ (.I(_0108_),
    .Z(_0109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0606_ (.A1(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .A2(_0109_),
    .ZN(_0110_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0607_ (.A1(_0106_),
    .A2(_0109_),
    .B(_0110_),
    .ZN(_0094_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0608_ (.I(net6),
    .ZN(_0111_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0609_ (.A1(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .A2(_0109_),
    .ZN(_0112_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0610_ (.A1(_0111_),
    .A2(_0109_),
    .B(_0112_),
    .ZN(_0093_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0611_ (.I(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .ZN(_0113_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0612_ (.A1(net5),
    .A2(_0108_),
    .ZN(_0114_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0613_ (.A1(_0113_),
    .A2(_0109_),
    .B(_0114_),
    .ZN(_0092_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0614_ (.I(net27),
    .ZN(_0115_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0615_ (.A1(\manchester_baby_instance.CIRCUIT_0.IR.q[4] ),
    .A2(_0109_),
    .ZN(_0116_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0616_ (.A1(_0115_),
    .A2(_0109_),
    .B(_0116_),
    .ZN(_0091_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _0617_ (.I(net26),
    .Z(_0117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0618_ (.I0(_0117_),
    .I1(\manchester_baby_instance.CIRCUIT_0.IR.q[3] ),
    .S(_0108_),
    .Z(_0118_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0619_ (.I(_0118_),
    .Z(_0090_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _0620_ (.I(net23),
    .Z(_0119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0621_ (.I0(_0119_),
    .I1(\manchester_baby_instance.CIRCUIT_0.IR.q[2] ),
    .S(_0108_),
    .Z(_0120_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0622_ (.I(_0120_),
    .Z(_0089_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0623_ (.I(net12),
    .ZN(_0121_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0624_ (.A1(\manchester_baby_instance.CIRCUIT_0.IR.q[1] ),
    .A2(_0109_),
    .ZN(_0122_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0625_ (.A1(_0121_),
    .A2(_0109_),
    .B(_0122_),
    .ZN(_0088_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0626_ (.I(net1),
    .ZN(_0123_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0627_ (.A1(\manchester_baby_instance.CIRCUIT_0.IR.q[0] ),
    .A2(_0108_),
    .ZN(_0124_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0628_ (.A1(_0123_),
    .A2(_0109_),
    .B(_0124_),
    .ZN(_0087_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0629_ (.I(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .ZN(_0125_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _0630_ (.A1(_0125_),
    .A2(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .A3(_0102_),
    .Z(_0126_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0631_ (.I(net24),
    .ZN(_0127_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0632_ (.A1(net63),
    .A2(_0127_),
    .ZN(_0128_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0633_ (.I(net16),
    .ZN(_0129_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0634_ (.A1(net55),
    .A2(_0129_),
    .ZN(_0130_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0635_ (.I(net54),
    .ZN(_0131_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0636_ (.A1(_0131_),
    .A2(net15),
    .ZN(_0132_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0637_ (.I(net53),
    .ZN(_0133_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0638_ (.A1(_0133_),
    .A2(net14),
    .Z(_0134_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0639_ (.A1(net52),
    .A2(net13),
    .Z(_0135_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0640_ (.I(_0135_),
    .ZN(_0136_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0641_ (.A1(_0134_),
    .A2(_0136_),
    .ZN(_0137_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0642_ (.I(net49),
    .ZN(_0138_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0643_ (.A1(_0138_),
    .A2(net10),
    .ZN(_0139_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _0644_ (.I(net11),
    .ZN(_0140_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0645_ (.A1(net50),
    .A2(_0140_),
    .Z(_0141_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0646_ (.A1(net49),
    .A2(net10),
    .Z(_0142_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0647_ (.A1(net50),
    .A2(net11),
    .Z(_0143_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0648_ (.A1(_0142_),
    .A2(_0143_),
    .ZN(_0144_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0649_ (.I(net9),
    .ZN(_0145_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0650_ (.A1(net48),
    .A2(_0145_),
    .ZN(_0146_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0651_ (.I(net8),
    .ZN(_0147_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0652_ (.A1(net47),
    .A2(_0147_),
    .ZN(_0148_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0653_ (.A1(net48),
    .A2(_0145_),
    .ZN(_0149_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0654_ (.A1(_0146_),
    .A2(_0148_),
    .B(_0149_),
    .ZN(_0150_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0655_ (.A1(net50),
    .A2(_0140_),
    .ZN(_0151_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0656_ (.I(_0151_),
    .ZN(_0152_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _0657_ (.A1(_0139_),
    .A2(_0141_),
    .B1(_0144_),
    .B2(_0150_),
    .C(_0152_),
    .ZN(_0153_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0658_ (.A1(_0133_),
    .A2(net14),
    .ZN(_0154_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0659_ (.I(net52),
    .ZN(_0155_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0660_ (.A1(_0155_),
    .A2(net13),
    .ZN(_0156_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0661_ (.A1(_0133_),
    .A2(net14),
    .ZN(_0157_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0662_ (.A1(_0154_),
    .A2(_0156_),
    .B(_0157_),
    .ZN(_0158_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0663_ (.A1(_0137_),
    .A2(_0153_),
    .B(_0158_),
    .ZN(_0159_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0664_ (.A1(_0131_),
    .A2(net15),
    .ZN(_0160_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0665_ (.A1(net55),
    .A2(_0129_),
    .B1(_0132_),
    .B2(_0159_),
    .C(_0160_),
    .ZN(_0161_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0666_ (.A1(_0130_),
    .A2(_0161_),
    .ZN(_0162_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0667_ (.A1(net7),
    .A2(net46),
    .Z(_0163_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0668_ (.A1(_0111_),
    .A2(net45),
    .Z(_0164_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0669_ (.I(_0164_),
    .ZN(_0165_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0670_ (.A1(net5),
    .A2(net44),
    .Z(_0166_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0671_ (.A1(net43),
    .A2(net4),
    .Z(_0167_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0672_ (.A1(_0163_),
    .A2(_0165_),
    .A3(_0166_),
    .A4(_0167_),
    .ZN(_0168_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0673_ (.I(net3),
    .ZN(_0169_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0674_ (.A1(net41),
    .A2(net2),
    .Z(_0170_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0675_ (.A1(net42),
    .A2(net3),
    .Z(_0171_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0676_ (.A1(_0170_),
    .A2(_0171_),
    .ZN(_0172_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0677_ (.I(net71),
    .ZN(_0173_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0678_ (.I(net31),
    .ZN(_0174_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0679_ (.I(net32),
    .ZN(_0175_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0680_ (.A1(net70),
    .A2(_0174_),
    .B1(_0175_),
    .B2(net71),
    .ZN(_0176_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0681_ (.A1(_0173_),
    .A2(net32),
    .B(_0176_),
    .ZN(_0177_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0682_ (.I(net42),
    .ZN(_0178_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0683_ (.I(net41),
    .ZN(_0179_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0684_ (.A1(_0178_),
    .A2(net3),
    .B(net2),
    .C(_0179_),
    .ZN(_0180_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0685_ (.A1(net42),
    .A2(_0169_),
    .B1(_0172_),
    .B2(_0177_),
    .C(_0180_),
    .ZN(_0181_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0686_ (.I(_0181_),
    .ZN(_0182_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0687_ (.I(net30),
    .ZN(_0183_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0688_ (.A1(net69),
    .A2(_0183_),
    .Z(_0184_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0689_ (.I(net29),
    .ZN(_0185_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0690_ (.A1(net68),
    .A2(_0185_),
    .Z(_0186_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0691_ (.A1(_0184_),
    .A2(_0186_),
    .ZN(_0187_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0692_ (.A1(net67),
    .A2(net28),
    .Z(_0188_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0693_ (.I(net65),
    .ZN(_0189_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0694_ (.A1(_0117_),
    .A2(_0189_),
    .ZN(_0190_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0695_ (.I(net62),
    .ZN(_0191_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _0696_ (.A1(_0117_),
    .A2(_0189_),
    .B(_0191_),
    .C(_0119_),
    .ZN(_0192_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0697_ (.A1(_0121_),
    .A2(net51),
    .ZN(_0193_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0698_ (.A1(net12),
    .A2(net51),
    .ZN(_0194_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0699_ (.A1(_0123_),
    .A2(net40),
    .B(_0194_),
    .ZN(_0195_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0700_ (.A1(_0119_),
    .A2(net62),
    .ZN(_0196_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0701_ (.A1(_0117_),
    .A2(net65),
    .ZN(_0197_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0702_ (.A1(_0196_),
    .A2(_0197_),
    .ZN(_0198_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0703_ (.A1(_0193_),
    .A2(_0195_),
    .B(_0198_),
    .ZN(_0199_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0704_ (.A1(net27),
    .A2(net66),
    .Z(_0200_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0705_ (.I(_0200_),
    .ZN(_0201_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _0706_ (.A1(_0190_),
    .A2(_0192_),
    .A3(_0199_),
    .B(_0201_),
    .ZN(_0202_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0707_ (.A1(_0184_),
    .A2(_0186_),
    .Z(_0203_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0708_ (.I(net28),
    .ZN(_0204_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0709_ (.A1(net67),
    .A2(_0204_),
    .ZN(_0205_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0710_ (.A1(_0115_),
    .A2(net66),
    .ZN(_0206_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0711_ (.A1(net67),
    .A2(_0204_),
    .ZN(_0207_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0712_ (.A1(_0205_),
    .A2(_0206_),
    .B(_0207_),
    .ZN(_0208_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0713_ (.A1(net69),
    .A2(_0183_),
    .ZN(_0209_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0714_ (.A1(net68),
    .A2(_0185_),
    .ZN(_0210_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0715_ (.A1(_0209_),
    .A2(_0210_),
    .ZN(_0211_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0716_ (.A1(net69),
    .A2(_0183_),
    .B1(_0203_),
    .B2(_0208_),
    .C(_0211_),
    .ZN(_0212_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _0717_ (.A1(_0187_),
    .A2(_0188_),
    .A3(_0202_),
    .B(_0212_),
    .ZN(_0213_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0718_ (.A1(_0173_),
    .A2(net32),
    .Z(_0214_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0719_ (.A1(net70),
    .A2(_0174_),
    .Z(_0215_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0720_ (.A1(_0214_),
    .A2(_0215_),
    .Z(_0216_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0721_ (.A1(_0172_),
    .A2(_0216_),
    .Z(_0217_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0722_ (.A1(_0168_),
    .A2(_0217_),
    .Z(_0218_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0723_ (.A1(_0168_),
    .A2(_0182_),
    .B1(_0213_),
    .B2(_0218_),
    .ZN(_0219_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0724_ (.A1(_0163_),
    .A2(_0165_),
    .ZN(_0220_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0725_ (.I(net44),
    .ZN(_0221_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0726_ (.A1(net5),
    .A2(_0221_),
    .ZN(_0222_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0727_ (.I(net43),
    .ZN(_0223_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0728_ (.A1(_0223_),
    .A2(net4),
    .ZN(_0224_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0729_ (.A1(net5),
    .A2(_0221_),
    .ZN(_0225_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0730_ (.A1(_0222_),
    .A2(_0224_),
    .B(_0225_),
    .ZN(_0226_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0731_ (.I(_0226_),
    .ZN(_0227_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0732_ (.A1(_0106_),
    .A2(net46),
    .ZN(_0228_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0733_ (.A1(_0111_),
    .A2(net45),
    .ZN(_0229_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0734_ (.A1(_0228_),
    .A2(_0229_),
    .ZN(_0230_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0735_ (.A1(_0106_),
    .A2(net46),
    .B1(_0220_),
    .B2(_0227_),
    .C(_0230_),
    .ZN(_0231_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0736_ (.A1(net48),
    .A2(net9),
    .Z(_0232_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0737_ (.A1(net47),
    .A2(_0147_),
    .Z(_0233_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0738_ (.I(_0233_),
    .ZN(_0234_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0739_ (.A1(_0232_),
    .A2(_0234_),
    .ZN(_0235_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0740_ (.A1(_0144_),
    .A2(_0235_),
    .ZN(_0236_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0741_ (.A1(net55),
    .A2(net16),
    .Z(_0237_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0742_ (.A1(net54),
    .A2(net15),
    .Z(_0238_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0743_ (.A1(_0137_),
    .A2(_0236_),
    .A3(_0237_),
    .A4(_0238_),
    .Z(_0239_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0744_ (.A1(_0219_),
    .A2(_0231_),
    .B(_0239_),
    .ZN(_0240_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0745_ (.A1(net59),
    .A2(net20),
    .Z(_0241_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0746_ (.I(_0241_),
    .ZN(_0242_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0747_ (.I(net19),
    .ZN(_0243_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0748_ (.A1(net58),
    .A2(_0243_),
    .Z(_0244_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0749_ (.A1(_0242_),
    .A2(_0244_),
    .ZN(_0245_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0750_ (.I(net57),
    .ZN(_0246_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0751_ (.A1(_0246_),
    .A2(net18),
    .Z(_0247_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0752_ (.A1(net56),
    .A2(net17),
    .Z(_0248_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0753_ (.I(_0248_),
    .ZN(_0249_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0754_ (.A1(_0247_),
    .A2(_0249_),
    .ZN(_0250_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0755_ (.A1(_0245_),
    .A2(_0250_),
    .ZN(_0251_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0756_ (.A1(_0162_),
    .A2(_0240_),
    .B(_0251_),
    .ZN(_0252_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0757_ (.I(net59),
    .ZN(_0253_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0758_ (.A1(_0253_),
    .A2(net20),
    .ZN(_0254_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0759_ (.A1(net58),
    .A2(_0243_),
    .ZN(_0255_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0760_ (.I(_0255_),
    .ZN(_0256_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0761_ (.A1(_0246_),
    .A2(net18),
    .ZN(_0257_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0762_ (.I(net17),
    .ZN(_0258_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0763_ (.A1(net56),
    .A2(_0258_),
    .ZN(_0259_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0764_ (.A1(_0246_),
    .A2(net18),
    .B(_0259_),
    .ZN(_0260_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0765_ (.A1(_0257_),
    .A2(_0260_),
    .ZN(_0261_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0766_ (.A1(_0253_),
    .A2(net20),
    .B1(_0245_),
    .B2(_0261_),
    .ZN(_0262_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0767_ (.A1(_0254_),
    .A2(_0256_),
    .B(_0262_),
    .ZN(_0263_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0768_ (.I(net22),
    .ZN(_0264_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0769_ (.A1(net61),
    .A2(_0264_),
    .Z(_0265_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0770_ (.I(net60),
    .ZN(_0266_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0771_ (.A1(_0266_),
    .A2(net21),
    .Z(_0267_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0772_ (.A1(_0265_),
    .A2(_0267_),
    .ZN(_0268_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0773_ (.A1(_0252_),
    .A2(_0263_),
    .B(_0268_),
    .ZN(_0269_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0774_ (.A1(net61),
    .A2(_0264_),
    .ZN(_0270_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0775_ (.A1(_0266_),
    .A2(net21),
    .ZN(_0271_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0776_ (.A1(net61),
    .A2(_0264_),
    .B(_0271_),
    .ZN(_0272_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0777_ (.A1(_0270_),
    .A2(_0272_),
    .ZN(_0273_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0778_ (.A1(net63),
    .A2(_0127_),
    .Z(_0274_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0779_ (.A1(_0269_),
    .A2(_0273_),
    .B(_0274_),
    .ZN(_0275_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0780_ (.A1(net64),
    .A2(net25),
    .Z(_0276_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0781_ (.A1(_0128_),
    .A2(_0275_),
    .A3(_0276_),
    .Z(_0277_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0782_ (.A1(_0128_),
    .A2(_0275_),
    .B(_0276_),
    .ZN(_0278_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0783_ (.A1(_0125_),
    .A2(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .ZN(_0279_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _0784_ (.A1(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .A2(_0102_),
    .A3(_0279_),
    .Z(_0280_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0785_ (.I(_0280_),
    .Z(_0281_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0786_ (.I(net20),
    .ZN(_0282_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0787_ (.I(net10),
    .ZN(_0283_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0788_ (.A1(_0117_),
    .A2(net23),
    .A3(net12),
    .A4(net1),
    .Z(_0284_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0789_ (.A1(net27),
    .A2(net28),
    .Z(_0285_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0790_ (.A1(net29),
    .A2(net30),
    .A3(_0284_),
    .A4(_0285_),
    .Z(_0286_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0791_ (.A1(net31),
    .A2(net32),
    .A3(net2),
    .A4(_0286_),
    .ZN(_0287_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0792_ (.A1(net5),
    .A2(net4),
    .ZN(_0288_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0793_ (.A1(net7),
    .A2(net6),
    .ZN(_0289_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0794_ (.A1(_0169_),
    .A2(_0287_),
    .A3(_0288_),
    .A4(_0289_),
    .Z(_0290_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _0795_ (.A1(_0147_),
    .A2(_0145_),
    .A3(_0283_),
    .A4(_0290_),
    .Z(_0291_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0796_ (.A1(net13),
    .A2(net14),
    .ZN(_0292_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0797_ (.A1(net15),
    .A2(net16),
    .ZN(_0293_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0798_ (.A1(_0140_),
    .A2(_0291_),
    .A3(_0292_),
    .A4(_0293_),
    .ZN(_0294_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _0799_ (.A1(net17),
    .A2(net18),
    .A3(_0294_),
    .Z(_0295_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0800_ (.A1(net19),
    .A2(_0295_),
    .ZN(_0296_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0801_ (.A1(_0282_),
    .A2(_0296_),
    .ZN(_0297_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0802_ (.A1(net21),
    .A2(net22),
    .A3(net24),
    .A4(_0297_),
    .ZN(_0298_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0803_ (.A1(net25),
    .A2(_0298_),
    .Z(_0299_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0804_ (.A1(_0126_),
    .A2(_0277_),
    .A3(_0278_),
    .B1(_0281_),
    .B2(_0299_),
    .ZN(_0300_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0805_ (.A1(_0125_),
    .A2(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .A3(_0102_),
    .ZN(_0301_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0806_ (.A1(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .A2(_0102_),
    .A3(_0279_),
    .ZN(_0302_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0807_ (.A1(_0301_),
    .A2(_0302_),
    .B(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .ZN(_0303_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _0808_ (.I(_0303_),
    .Z(_0304_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0809_ (.I0(_0300_),
    .I1(net64),
    .S(_0304_),
    .Z(_0305_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0810_ (.I(_0305_),
    .Z(_0086_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0811_ (.A1(net21),
    .A2(_0297_),
    .ZN(_0306_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0812_ (.A1(_0264_),
    .A2(_0306_),
    .B(_0127_),
    .ZN(_0307_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0813_ (.A1(_0301_),
    .A2(_0275_),
    .ZN(_0308_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0814_ (.A1(_0274_),
    .A2(_0269_),
    .A3(_0273_),
    .ZN(_0309_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0815_ (.A1(_0281_),
    .A2(_0298_),
    .A3(_0307_),
    .B1(_0308_),
    .B2(_0309_),
    .ZN(_0310_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0816_ (.I0(_0310_),
    .I1(net63),
    .S(_0304_),
    .Z(_0311_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0817_ (.I(_0311_),
    .Z(_0085_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _0818_ (.I(_0303_),
    .Z(_0312_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0819_ (.I(_0312_),
    .Z(_0313_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0820_ (.I(_0302_),
    .Z(_0314_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0821_ (.A1(_0264_),
    .A2(_0306_),
    .Z(_0315_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0822_ (.A1(_0252_),
    .A2(_0263_),
    .ZN(_0316_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0823_ (.A1(_0316_),
    .A2(_0267_),
    .B(_0271_),
    .ZN(_0317_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0824_ (.A1(_0265_),
    .A2(_0317_),
    .ZN(_0318_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _0825_ (.I(_0301_),
    .Z(_0319_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0826_ (.A1(_0314_),
    .A2(_0315_),
    .B1(_0318_),
    .B2(_0319_),
    .ZN(_0320_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _0827_ (.I(_0312_),
    .Z(_0321_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0828_ (.A1(net61),
    .A2(_0321_),
    .ZN(_0322_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0829_ (.A1(_0313_),
    .A2(_0320_),
    .B(_0322_),
    .ZN(_0084_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0830_ (.I(_0301_),
    .Z(_0323_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0831_ (.A1(_0316_),
    .A2(_0267_),
    .Z(_0324_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0832_ (.A1(net21),
    .A2(_0297_),
    .Z(_0325_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0833_ (.A1(_0323_),
    .A2(_0324_),
    .B1(_0325_),
    .B2(_0314_),
    .ZN(_0326_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0834_ (.A1(net60),
    .A2(_0321_),
    .ZN(_0327_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0835_ (.A1(_0313_),
    .A2(_0326_),
    .B(_0327_),
    .ZN(_0083_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0836_ (.A1(net20),
    .A2(_0296_),
    .Z(_0328_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0837_ (.A1(_0162_),
    .A2(_0240_),
    .ZN(_0329_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0838_ (.A1(_0329_),
    .A2(_0250_),
    .B(_0261_),
    .ZN(_0330_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0839_ (.A1(_0244_),
    .A2(_0330_),
    .B(_0256_),
    .ZN(_0331_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0840_ (.A1(_0242_),
    .A2(_0331_),
    .Z(_0332_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0841_ (.A1(_0281_),
    .A2(_0328_),
    .B1(_0332_),
    .B2(_0126_),
    .ZN(_0333_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0842_ (.I0(_0333_),
    .I1(net59),
    .S(_0304_),
    .Z(_0334_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0843_ (.I(_0334_),
    .Z(_0082_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0844_ (.A1(_0244_),
    .A2(_0330_),
    .Z(_0335_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0845_ (.A1(net19),
    .A2(_0295_),
    .Z(_0336_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0846_ (.A1(_0323_),
    .A2(_0335_),
    .B1(_0336_),
    .B2(_0314_),
    .ZN(_0337_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0847_ (.A1(net58),
    .A2(_0321_),
    .ZN(_0338_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0848_ (.A1(_0313_),
    .A2(_0337_),
    .B(_0338_),
    .ZN(_0081_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0849_ (.A1(net17),
    .A2(_0294_),
    .B(net18),
    .ZN(_0339_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0850_ (.A1(_0295_),
    .A2(_0339_),
    .Z(_0340_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0851_ (.A1(_0329_),
    .A2(_0248_),
    .B(_0259_),
    .ZN(_0341_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0852_ (.A1(_0247_),
    .A2(_0341_),
    .Z(_0342_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0853_ (.A1(_0314_),
    .A2(_0340_),
    .B1(_0342_),
    .B2(_0319_),
    .ZN(_0343_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0854_ (.A1(net57),
    .A2(_0321_),
    .ZN(_0344_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0855_ (.A1(_0313_),
    .A2(_0343_),
    .B(_0344_),
    .ZN(_0080_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0856_ (.A1(net17),
    .A2(_0294_),
    .Z(_0345_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0857_ (.A1(_0329_),
    .A2(_0248_),
    .Z(_0346_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0858_ (.A1(_0314_),
    .A2(_0345_),
    .B1(_0346_),
    .B2(_0319_),
    .ZN(_0347_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0859_ (.A1(net56),
    .A2(_0321_),
    .ZN(_0348_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0860_ (.A1(_0313_),
    .A2(_0347_),
    .B(_0348_),
    .ZN(_0079_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0861_ (.A1(_0140_),
    .A2(_0291_),
    .A3(_0292_),
    .ZN(_0349_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0862_ (.A1(net15),
    .A2(_0349_),
    .B(net16),
    .ZN(_0350_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0863_ (.A1(_0294_),
    .A2(_0350_),
    .Z(_0351_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0864_ (.A1(_0219_),
    .A2(_0231_),
    .ZN(_0352_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0865_ (.I(_0236_),
    .ZN(_0353_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0866_ (.A1(_0144_),
    .A2(_0150_),
    .ZN(_0354_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0867_ (.A1(_0151_),
    .A2(_0354_),
    .ZN(_0355_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0868_ (.A1(_0139_),
    .A2(_0141_),
    .B1(_0352_),
    .B2(_0353_),
    .C(_0355_),
    .ZN(_0356_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0869_ (.A1(_0137_),
    .A2(_0356_),
    .B(_0158_),
    .ZN(_0357_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0870_ (.A1(_0132_),
    .A2(_0357_),
    .B(_0160_),
    .ZN(_0358_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0871_ (.A1(_0237_),
    .A2(_0358_),
    .Z(_0359_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0872_ (.A1(_0314_),
    .A2(_0351_),
    .B1(_0359_),
    .B2(_0319_),
    .ZN(_0360_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0873_ (.I(_0303_),
    .Z(_0361_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0874_ (.A1(net55),
    .A2(_0361_),
    .ZN(_0362_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0875_ (.A1(_0313_),
    .A2(_0360_),
    .B(_0362_),
    .ZN(_0078_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0876_ (.A1(net15),
    .A2(_0349_),
    .ZN(_0363_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0877_ (.A1(_0238_),
    .A2(_0357_),
    .Z(_0364_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0878_ (.A1(_0281_),
    .A2(_0363_),
    .B1(_0364_),
    .B2(_0126_),
    .ZN(_0365_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0879_ (.I0(_0365_),
    .I1(net54),
    .S(_0312_),
    .Z(_0366_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0880_ (.I(_0366_),
    .Z(_0077_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0881_ (.A1(_0135_),
    .A2(_0356_),
    .ZN(_0367_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0882_ (.A1(_0156_),
    .A2(_0367_),
    .ZN(_0368_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0883_ (.A1(_0134_),
    .A2(_0368_),
    .Z(_0369_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0884_ (.A1(_0140_),
    .A2(_0291_),
    .ZN(_0370_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0885_ (.A1(net13),
    .A2(_0370_),
    .B(net14),
    .ZN(_0371_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0886_ (.A1(_0302_),
    .A2(_0349_),
    .A3(_0371_),
    .ZN(_0372_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0887_ (.A1(_0126_),
    .A2(_0369_),
    .B(_0372_),
    .ZN(_0373_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0888_ (.I0(_0373_),
    .I1(net53),
    .S(_0312_),
    .Z(_0374_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0889_ (.I(_0374_),
    .Z(_0076_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0890_ (.A1(net13),
    .A2(_0370_),
    .Z(_0375_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0891_ (.A1(_0135_),
    .A2(_0356_),
    .ZN(_0376_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0892_ (.A1(_0126_),
    .A2(_0367_),
    .ZN(_0377_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0893_ (.A1(_0314_),
    .A2(_0375_),
    .B1(_0376_),
    .B2(_0377_),
    .ZN(_0378_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0894_ (.A1(net52),
    .A2(_0361_),
    .ZN(_0379_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0895_ (.A1(_0313_),
    .A2(_0378_),
    .B(_0379_),
    .ZN(_0075_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _0896_ (.I(_0302_),
    .Z(_0380_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0897_ (.A1(_0140_),
    .A2(_0291_),
    .Z(_0381_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0898_ (.A1(_0352_),
    .A2(_0235_),
    .B(_0150_),
    .ZN(_0382_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0899_ (.A1(_0142_),
    .A2(_0382_),
    .Z(_0383_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0900_ (.A1(_0138_),
    .A2(net10),
    .B(_0383_),
    .ZN(_0384_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0901_ (.A1(_0143_),
    .A2(_0384_),
    .ZN(_0385_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0902_ (.A1(_0380_),
    .A2(_0381_),
    .B1(_0385_),
    .B2(_0319_),
    .ZN(_0386_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0903_ (.A1(net50),
    .A2(_0361_),
    .ZN(_0387_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0904_ (.A1(_0313_),
    .A2(_0386_),
    .B(_0387_),
    .ZN(_0074_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0905_ (.I(_0312_),
    .Z(_0388_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0906_ (.A1(_0147_),
    .A2(_0290_),
    .ZN(_0389_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0907_ (.A1(net9),
    .A2(_0389_),
    .ZN(_0390_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0908_ (.A1(_0283_),
    .A2(_0390_),
    .Z(_0391_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0909_ (.A1(_0301_),
    .A2(_0383_),
    .ZN(_0392_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0910_ (.A1(_0142_),
    .A2(_0382_),
    .B(_0392_),
    .ZN(_0393_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0911_ (.A1(_0314_),
    .A2(_0391_),
    .B(_0393_),
    .ZN(_0394_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0912_ (.A1(net49),
    .A2(_0361_),
    .ZN(_0395_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0913_ (.A1(_0388_),
    .A2(_0394_),
    .B(_0395_),
    .ZN(_0073_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0914_ (.A1(net9),
    .A2(_0389_),
    .Z(_0396_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0915_ (.A1(_0352_),
    .A2(_0233_),
    .ZN(_0397_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0916_ (.A1(_0148_),
    .A2(_0397_),
    .ZN(_0398_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0917_ (.A1(_0232_),
    .A2(_0398_),
    .ZN(_0399_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0918_ (.A1(_0380_),
    .A2(_0396_),
    .B1(_0399_),
    .B2(_0319_),
    .ZN(_0400_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0919_ (.A1(net48),
    .A2(_0361_),
    .ZN(_0401_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0920_ (.A1(_0388_),
    .A2(_0400_),
    .B(_0401_),
    .ZN(_0072_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0921_ (.A1(_0352_),
    .A2(_0233_),
    .Z(_0402_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0922_ (.A1(_0147_),
    .A2(_0290_),
    .Z(_0403_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0923_ (.A1(_0323_),
    .A2(_0402_),
    .B1(_0403_),
    .B2(_0314_),
    .ZN(_0404_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0924_ (.A1(net47),
    .A2(_0361_),
    .ZN(_0405_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0925_ (.A1(_0388_),
    .A2(_0404_),
    .B(_0405_),
    .ZN(_0071_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0926_ (.A1(_0213_),
    .A2(_0217_),
    .B(_0182_),
    .ZN(_0406_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _0927_ (.A1(_0166_),
    .A2(_0167_),
    .A3(_0406_),
    .B(_0226_),
    .ZN(_0407_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0928_ (.A1(_0164_),
    .A2(_0407_),
    .ZN(_0408_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0929_ (.A1(_0229_),
    .A2(_0408_),
    .ZN(_0409_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0930_ (.A1(_0163_),
    .A2(_0409_),
    .ZN(_0410_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0931_ (.A1(_0169_),
    .A2(_0287_),
    .A3(_0288_),
    .ZN(_0411_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0932_ (.A1(net6),
    .A2(_0411_),
    .B(net7),
    .ZN(_0412_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0933_ (.A1(_0281_),
    .A2(_0290_),
    .ZN(_0413_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0934_ (.A1(_0323_),
    .A2(_0410_),
    .B1(_0412_),
    .B2(_0413_),
    .ZN(_0414_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0935_ (.A1(net46),
    .A2(_0361_),
    .ZN(_0415_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0936_ (.A1(_0388_),
    .A2(_0414_),
    .B(_0415_),
    .ZN(_0070_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0937_ (.A1(net6),
    .A2(_0411_),
    .Z(_0416_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0938_ (.A1(_0164_),
    .A2(_0407_),
    .Z(_0417_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0939_ (.A1(_0380_),
    .A2(_0416_),
    .B1(_0417_),
    .B2(_0319_),
    .ZN(_0418_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0940_ (.A1(net45),
    .A2(_0361_),
    .ZN(_0419_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0941_ (.A1(_0388_),
    .A2(_0418_),
    .B(_0419_),
    .ZN(_0069_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0942_ (.A1(_0169_),
    .A2(_0287_),
    .ZN(_0420_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0943_ (.A1(net4),
    .A2(_0420_),
    .B(net5),
    .ZN(_0421_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0944_ (.A1(_0411_),
    .A2(_0421_),
    .Z(_0422_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0945_ (.A1(_0167_),
    .A2(_0406_),
    .ZN(_0423_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0946_ (.A1(_0224_),
    .A2(_0423_),
    .ZN(_0424_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0947_ (.A1(_0166_),
    .A2(_0424_),
    .Z(_0425_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0948_ (.A1(_0380_),
    .A2(_0422_),
    .B1(_0425_),
    .B2(_0319_),
    .ZN(_0426_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0949_ (.A1(net44),
    .A2(_0361_),
    .ZN(_0427_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0950_ (.A1(_0388_),
    .A2(_0426_),
    .B(_0427_),
    .ZN(_0068_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0951_ (.A1(net4),
    .A2(_0420_),
    .Z(_0428_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0952_ (.A1(_0167_),
    .A2(_0406_),
    .ZN(_0429_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0953_ (.A1(_0126_),
    .A2(_0423_),
    .ZN(_0430_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0954_ (.A1(_0380_),
    .A2(_0428_),
    .B1(_0429_),
    .B2(_0430_),
    .ZN(_0431_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0955_ (.A1(net43),
    .A2(_0361_),
    .ZN(_0432_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0956_ (.A1(_0388_),
    .A2(_0431_),
    .B(_0432_),
    .ZN(_0067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0957_ (.A1(_0169_),
    .A2(_0287_),
    .Z(_0433_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0958_ (.A1(_0179_),
    .A2(net2),
    .ZN(_0434_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0959_ (.A1(_0213_),
    .A2(_0216_),
    .B(_0177_),
    .ZN(_0435_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0960_ (.A1(_0170_),
    .A2(_0435_),
    .ZN(_0436_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0961_ (.A1(_0434_),
    .A2(_0436_),
    .ZN(_0437_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0962_ (.A1(_0171_),
    .A2(_0437_),
    .Z(_0438_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0963_ (.A1(_0380_),
    .A2(_0433_),
    .B1(_0438_),
    .B2(_0319_),
    .ZN(_0439_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0964_ (.A1(net42),
    .A2(_0304_),
    .ZN(_0440_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0965_ (.A1(_0388_),
    .A2(_0439_),
    .B(_0440_),
    .ZN(_0066_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0966_ (.A1(net31),
    .A2(net32),
    .A3(_0286_),
    .B(net2),
    .ZN(_0441_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0967_ (.A1(_0281_),
    .A2(_0287_),
    .ZN(_0442_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0968_ (.A1(_0170_),
    .A2(_0435_),
    .ZN(_0443_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0969_ (.A1(_0126_),
    .A2(_0436_),
    .ZN(_0444_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0970_ (.A1(_0441_),
    .A2(_0442_),
    .B1(_0443_),
    .B2(_0444_),
    .ZN(_0445_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0971_ (.A1(net41),
    .A2(_0304_),
    .ZN(_0446_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0972_ (.A1(_0388_),
    .A2(_0445_),
    .B(_0446_),
    .ZN(_0065_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0973_ (.A1(net31),
    .A2(_0286_),
    .ZN(_0447_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0974_ (.A1(_0175_),
    .A2(_0447_),
    .Z(_0448_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0975_ (.A1(net70),
    .A2(_0174_),
    .ZN(_0449_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0976_ (.A1(_0213_),
    .A2(_0215_),
    .ZN(_0450_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0977_ (.A1(_0449_),
    .A2(_0450_),
    .ZN(_0451_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0978_ (.A1(_0214_),
    .A2(_0451_),
    .Z(_0452_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0979_ (.A1(_0380_),
    .A2(_0448_),
    .B1(_0452_),
    .B2(_0319_),
    .ZN(_0453_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0980_ (.A1(net71),
    .A2(_0304_),
    .ZN(_0454_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0981_ (.A1(_0388_),
    .A2(_0453_),
    .B(_0454_),
    .ZN(_0064_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0982_ (.A1(net31),
    .A2(_0286_),
    .ZN(_0455_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0983_ (.A1(_0281_),
    .A2(_0447_),
    .ZN(_0456_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0984_ (.A1(_0213_),
    .A2(_0215_),
    .Z(_0457_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0985_ (.A1(_0455_),
    .A2(_0456_),
    .B1(_0457_),
    .B2(_0323_),
    .ZN(_0458_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0986_ (.A1(net70),
    .A2(_0304_),
    .ZN(_0459_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0987_ (.A1(_0321_),
    .A2(_0458_),
    .B(_0459_),
    .ZN(_0063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0988_ (.A1(_0284_),
    .A2(_0285_),
    .Z(_0460_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0989_ (.A1(net29),
    .A2(_0460_),
    .ZN(_0461_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0990_ (.A1(_0183_),
    .A2(_0461_),
    .Z(_0462_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0991_ (.A1(_0188_),
    .A2(_0202_),
    .ZN(_0463_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0992_ (.A1(_0463_),
    .A2(_0208_),
    .B(_0186_),
    .ZN(_0464_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0993_ (.A1(_0210_),
    .A2(_0464_),
    .ZN(_0465_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0994_ (.A1(_0184_),
    .A2(_0465_),
    .Z(_0466_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0995_ (.A1(_0380_),
    .A2(_0462_),
    .B1(_0466_),
    .B2(_0323_),
    .ZN(_0467_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0996_ (.A1(net69),
    .A2(_0304_),
    .ZN(_0468_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0997_ (.A1(_0321_),
    .A2(_0467_),
    .B(_0468_),
    .ZN(_0062_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0998_ (.A1(net29),
    .A2(_0460_),
    .ZN(_0469_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0999_ (.A1(_0281_),
    .A2(_0461_),
    .ZN(_0470_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1000_ (.A1(_0186_),
    .A2(_0463_),
    .A3(_0208_),
    .Z(_0471_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1001_ (.A1(_0301_),
    .A2(_0464_),
    .Z(_0472_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1002_ (.A1(_0469_),
    .A2(_0470_),
    .B1(_0471_),
    .B2(_0472_),
    .ZN(_0473_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1003_ (.A1(net68),
    .A2(_0304_),
    .ZN(_0474_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1004_ (.A1(_0321_),
    .A2(_0473_),
    .B(_0474_),
    .ZN(_0061_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1005_ (.A1(_0206_),
    .A2(_0202_),
    .ZN(_0475_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1006_ (.A1(_0188_),
    .A2(_0475_),
    .Z(_0476_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1007_ (.A1(net27),
    .A2(_0284_),
    .B(net28),
    .ZN(_0477_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1008_ (.A1(_0302_),
    .A2(_0460_),
    .A3(_0477_),
    .ZN(_0478_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1009_ (.A1(_0126_),
    .A2(_0476_),
    .B(_0478_),
    .ZN(_0479_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1010_ (.I0(_0479_),
    .I1(net67),
    .S(_0312_),
    .Z(_0480_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1011_ (.I(_0480_),
    .Z(_0060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1012_ (.A1(_0190_),
    .A2(_0192_),
    .A3(_0199_),
    .A4(_0201_),
    .Z(_0481_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1013_ (.A1(_0301_),
    .A2(_0202_),
    .Z(_0482_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1014_ (.A1(net27),
    .A2(_0284_),
    .Z(_0483_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1015_ (.A1(_0481_),
    .A2(_0482_),
    .B1(_0483_),
    .B2(_0314_),
    .ZN(_0484_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1016_ (.A1(net66),
    .A2(_0304_),
    .ZN(_0485_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1017_ (.A1(_0321_),
    .A2(_0484_),
    .B(_0485_),
    .ZN(_0059_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1018_ (.A1(_0193_),
    .A2(_0195_),
    .ZN(_0486_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1019_ (.A1(_0486_),
    .A2(_0196_),
    .ZN(_0487_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1020_ (.A1(_0119_),
    .A2(_0191_),
    .B(_0487_),
    .ZN(_0488_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1021_ (.A1(_0488_),
    .A2(_0197_),
    .Z(_0489_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1022_ (.A1(_0119_),
    .A2(net12),
    .A3(net1),
    .Z(_0490_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1023_ (.A1(_0302_),
    .A2(_0284_),
    .ZN(_0491_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1024_ (.A1(_0117_),
    .A2(_0490_),
    .B(_0491_),
    .ZN(_0492_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1025_ (.A1(_0323_),
    .A2(_0489_),
    .B(_0492_),
    .C(_0312_),
    .ZN(_0493_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1026_ (.A1(_0189_),
    .A2(_0313_),
    .B(_0493_),
    .ZN(_0058_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1027_ (.A1(_0486_),
    .A2(_0196_),
    .Z(_0494_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1028_ (.A1(net12),
    .A2(net1),
    .B(_0119_),
    .ZN(_0495_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1029_ (.A1(_0490_),
    .A2(_0495_),
    .Z(_0496_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1030_ (.A1(_0323_),
    .A2(_0494_),
    .B1(_0496_),
    .B2(_0380_),
    .C(_0312_),
    .ZN(_0497_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1031_ (.A1(_0191_),
    .A2(_0313_),
    .B(_0497_),
    .ZN(_0057_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1032_ (.A1(_0121_),
    .A2(net1),
    .Z(_0498_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1033_ (.A1(_0123_),
    .A2(net40),
    .A3(_0194_),
    .ZN(_0499_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1034_ (.A1(_0323_),
    .A2(_0195_),
    .ZN(_0500_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1035_ (.A1(_0281_),
    .A2(_0498_),
    .B1(_0499_),
    .B2(_0500_),
    .ZN(_0501_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1036_ (.I0(_0501_),
    .I1(net51),
    .S(_0312_),
    .Z(_0502_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1037_ (.I(_0502_),
    .Z(_0056_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1038_ (.I(net40),
    .ZN(_0503_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1039_ (.A1(_0503_),
    .A2(_0380_),
    .ZN(_0504_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1040_ (.A1(_0123_),
    .A2(_0323_),
    .B(_0312_),
    .ZN(_0505_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1041_ (.A1(_0123_),
    .A2(_0321_),
    .A3(_0504_),
    .B1(_0505_),
    .B2(_0503_),
    .ZN(_0055_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _1042_ (.A1(_0107_),
    .A2(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .A3(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ),
    .Z(_0506_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1043_ (.A1(_0107_),
    .A2(_0101_),
    .ZN(_0507_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1044_ (.A1(_0506_),
    .A2(_0507_),
    .ZN(_0508_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1045_ (.A1(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .A2(_0508_),
    .ZN(_0509_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1046_ (.A1(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .A2(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .Z(_0510_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1047_ (.A1(_0113_),
    .A2(_0506_),
    .A3(_0510_),
    .ZN(_0511_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1048_ (.A1(_0117_),
    .A2(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .ZN(_0512_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1049_ (.A1(_0119_),
    .A2(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .ZN(_0513_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1050_ (.I(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .Z(_0514_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1051_ (.A1(net12),
    .A2(_0514_),
    .ZN(_0515_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1052_ (.A1(net12),
    .A2(_0514_),
    .Z(_0516_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1053_ (.A1(net1),
    .A2(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .A3(_0516_),
    .ZN(_0517_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1054_ (.A1(_0515_),
    .A2(_0517_),
    .ZN(_0518_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1055_ (.A1(_0119_),
    .A2(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .B(_0518_),
    .ZN(_0519_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1056_ (.A1(_0513_),
    .A2(_0519_),
    .ZN(_0520_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1057_ (.A1(_0117_),
    .A2(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .B(_0520_),
    .ZN(_0521_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1058_ (.A1(_0512_),
    .A2(_0521_),
    .ZN(_0522_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1059_ (.A1(net27),
    .A2(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .A3(_0522_),
    .Z(_0523_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1060_ (.A1(_0511_),
    .A2(_0523_),
    .ZN(_0524_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1061_ (.A1(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .A2(_0103_),
    .A3(_0506_),
    .Z(_0525_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1062_ (.A1(_0507_),
    .A2(_0525_),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .ZN(_0526_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1063_ (.A1(net64),
    .A2(_0514_),
    .A3(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .Z(_0527_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1064_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A2(_0527_),
    .B(_0525_),
    .ZN(_0528_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1065_ (.A1(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .A2(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .A3(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .ZN(_0529_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1066_ (.I(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .Z(_0530_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1067_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A2(_0514_),
    .A3(_0530_),
    .ZN(_0531_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1068_ (.A1(_0529_),
    .A2(_0531_),
    .ZN(_0532_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1069_ (.I(_0532_),
    .ZN(_0533_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1070_ (.A1(_0526_),
    .A2(_0528_),
    .A3(_0533_),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .ZN(_0534_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1071_ (.A1(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .A2(_0506_),
    .A3(_0510_),
    .ZN(_0535_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1072_ (.A1(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .A2(_0103_),
    .A3(_0506_),
    .ZN(_0536_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1073_ (.A1(net64),
    .A2(_0536_),
    .ZN(_0537_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1074_ (.A1(_0507_),
    .A2(_0537_),
    .B(_0531_),
    .ZN(_0538_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1075_ (.I(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .ZN(_0539_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1076_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .A2(_0539_),
    .ZN(_0540_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1077_ (.A1(net27),
    .A2(_0535_),
    .B1(_0538_),
    .B2(_0540_),
    .ZN(_0541_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1078_ (.A1(_0524_),
    .A2(_0534_),
    .A3(_0541_),
    .Z(_0542_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1079_ (.A1(_0103_),
    .A2(_0510_),
    .ZN(_0543_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1080_ (.A1(_0506_),
    .A2(_0543_),
    .B(_0508_),
    .C(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .ZN(_0544_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1081_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .A2(_0544_),
    .ZN(_0545_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1082_ (.A1(_0509_),
    .A2(_0542_),
    .B(_0545_),
    .ZN(_0054_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1083_ (.A1(_0117_),
    .A2(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A3(_0520_),
    .Z(_0546_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1084_ (.A1(_0507_),
    .A2(_0537_),
    .B(_0531_),
    .C(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .ZN(_0547_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1085_ (.A1(_0117_),
    .A2(_0535_),
    .B1(_0546_),
    .B2(_0511_),
    .C(_0547_),
    .ZN(_0548_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1086_ (.A1(_0544_),
    .A2(_0528_),
    .A3(_0533_),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .ZN(_0549_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1087_ (.A1(_0509_),
    .A2(_0548_),
    .B(_0549_),
    .ZN(_0053_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1088_ (.A1(_0119_),
    .A2(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A3(_0518_),
    .Z(_0550_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1089_ (.A1(_0514_),
    .A2(_0530_),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .ZN(_0551_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1090_ (.A1(_0119_),
    .A2(_0535_),
    .ZN(_0552_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1091_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A2(_0527_),
    .B(_0528_),
    .ZN(_0553_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1092_ (.A1(_0532_),
    .A2(_0551_),
    .B(_0552_),
    .C(_0553_),
    .ZN(_0554_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1093_ (.A1(_0511_),
    .A2(_0550_),
    .B(_0554_),
    .ZN(_0555_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1094_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A2(_0544_),
    .ZN(_0556_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1095_ (.A1(_0509_),
    .A2(_0555_),
    .B(_0556_),
    .ZN(_0052_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1096_ (.A1(_0514_),
    .A2(_0530_),
    .Z(_0557_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1097_ (.A1(net64),
    .A2(_0530_),
    .B(_0514_),
    .ZN(_0558_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1098_ (.A1(net1),
    .A2(_0530_),
    .B(_0516_),
    .ZN(_0559_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1099_ (.A1(_0517_),
    .A2(_0511_),
    .ZN(_0560_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1100_ (.A1(_0525_),
    .A2(_0527_),
    .A3(_0558_),
    .B1(_0559_),
    .B2(_0560_),
    .ZN(_0561_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1101_ (.A1(net12),
    .A2(_0535_),
    .B1(_0557_),
    .B2(_0529_),
    .C(_0561_),
    .ZN(_0562_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1102_ (.A1(_0514_),
    .A2(_0544_),
    .ZN(_0563_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1103_ (.A1(_0509_),
    .A2(_0562_),
    .B(_0563_),
    .ZN(_0051_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1104_ (.A1(net64),
    .A2(_0530_),
    .Z(_0564_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1105_ (.A1(net1),
    .A2(_0530_),
    .Z(_0565_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1106_ (.A1(_0511_),
    .A2(_0565_),
    .ZN(_0566_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1107_ (.A1(_0530_),
    .A2(_0507_),
    .B(_0566_),
    .ZN(_0567_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1108_ (.A1(net1),
    .A2(_0535_),
    .B1(_0564_),
    .B2(_0536_),
    .C(_0567_),
    .ZN(_0568_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1109_ (.A1(_0530_),
    .A2(_0544_),
    .ZN(_0569_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1110_ (.A1(_0509_),
    .A2(_0568_),
    .B(_0569_),
    .ZN(_0050_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1111_ (.A1(\manchester_baby_instance.BASE_0.s_countReg[0] ),
    .A2(\manchester_baby_instance.BASE_0.s_countReg[1] ),
    .A3(\manchester_baby_instance.BASE_0.s_countReg[2] ),
    .ZN(\manchester_baby_instance.BASE_0.s_tickNext ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1112_ (.A1(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .A2(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .ZN(_0570_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1113_ (.A1(_0113_),
    .A2(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .A3(_0279_),
    .A4(_0570_),
    .ZN(_0571_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1114_ (.I(_0571_),
    .Z(net72),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1115_ (.A1(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .A2(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .Z(_0572_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1116_ (.I(_0572_),
    .Z(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1117_ (.A1(_0107_),
    .A2(_0570_),
    .Z(_0573_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1118_ (.I(_0573_),
    .Z(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1119_ (.A1(_0105_),
    .A2(net34),
    .Z(_0574_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1120_ (.I(_0574_),
    .Z(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1121_ (.A1(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .A2(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .A3(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ),
    .ZN(_0575_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _1122_ (.A1(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .A2(_0543_),
    .A3(_0570_),
    .B1(_0102_),
    .B2(_0510_),
    .ZN(_0576_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1123_ (.A1(_0530_),
    .A2(_0575_),
    .B1(_0576_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[0] ),
    .ZN(_0577_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1124_ (.I(_0577_),
    .ZN(net35),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1125_ (.A1(_0514_),
    .A2(_0575_),
    .B1(_0576_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[1] ),
    .ZN(_0578_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1126_ (.I(_0578_),
    .ZN(net36),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1127_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A2(_0575_),
    .B1(_0576_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[2] ),
    .ZN(_0579_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1128_ (.I(_0579_),
    .ZN(net37),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1129_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(_0575_),
    .B1(_0576_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[3] ),
    .ZN(_0580_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1130_ (.I(_0580_),
    .ZN(net38),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1131_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .A2(_0575_),
    .B1(_0576_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[4] ),
    .ZN(_0581_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1132_ (.I(_0581_),
    .ZN(net39),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1133_ (.I(\manchester_baby_instance.BASE_1.s_derivedClock ),
    .ZN(_0582_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1134_ (.A1(_0582_),
    .A2(\manchester_baby_instance.BASE_1.s_bufferRegs[0] ),
    .ZN(_0000_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1135_ (.I(net33),
    .Z(_0583_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1136_ (.I(_0583_),
    .Z(_0584_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1137_ (.I(_0584_),
    .Z(_0585_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1138_ (.I(_0585_),
    .ZN(_0001_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1139_ (.I(_0585_),
    .ZN(_0002_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1140_ (.I(_0585_),
    .ZN(_0003_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1141_ (.I(_0585_),
    .ZN(_0004_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1142_ (.I(_0585_),
    .ZN(_0005_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1143_ (.I(_0585_),
    .ZN(_0006_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1144_ (.I(_0585_),
    .ZN(_0007_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1145_ (.I(_0585_),
    .ZN(_0008_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1146_ (.I(_0585_),
    .ZN(_0009_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1147_ (.I(_0585_),
    .ZN(_0010_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1148_ (.I(_0583_),
    .Z(_0586_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1149_ (.I(_0586_),
    .ZN(_0011_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1150_ (.I(_0586_),
    .ZN(_0012_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1151_ (.I(_0586_),
    .ZN(_0013_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1152_ (.I(_0586_),
    .ZN(_0014_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1153_ (.I(_0586_),
    .ZN(_0015_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1154_ (.I(_0586_),
    .ZN(_0016_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1155_ (.I(_0586_),
    .ZN(_0017_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1156_ (.I(_0586_),
    .ZN(_0018_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1157_ (.I(_0586_),
    .ZN(_0019_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1158_ (.I(_0586_),
    .ZN(_0020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1159_ (.I(_0583_),
    .Z(_0587_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1160_ (.I(_0587_),
    .ZN(_0021_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1161_ (.I(_0587_),
    .ZN(_0022_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1162_ (.I(_0587_),
    .ZN(_0023_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1163_ (.I(_0587_),
    .ZN(_0024_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1164_ (.I(_0587_),
    .ZN(_0025_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1165_ (.I(_0587_),
    .ZN(_0026_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1166_ (.I(_0587_),
    .ZN(_0027_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1167_ (.I(_0587_),
    .ZN(_0028_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1168_ (.I(_0587_),
    .ZN(_0029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1169_ (.I(_0587_),
    .ZN(_0030_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1170_ (.I(_0583_),
    .Z(_0588_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1171_ (.I(_0588_),
    .ZN(_0031_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1172_ (.I(_0588_),
    .ZN(_0032_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1173_ (.I(_0588_),
    .ZN(_0033_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1174_ (.I(_0588_),
    .ZN(_0034_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1175_ (.I(_0588_),
    .ZN(_0035_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1176_ (.I(_0588_),
    .ZN(_0036_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1177_ (.I(_0588_),
    .ZN(_0037_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1178_ (.I(_0588_),
    .ZN(_0038_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1179_ (.I(_0588_),
    .ZN(_0039_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1180_ (.I(_0588_),
    .ZN(_0040_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1181_ (.I(_0584_),
    .ZN(_0041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1182_ (.I(_0584_),
    .ZN(_0042_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1183_ (.I(_0584_),
    .ZN(_0043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1184_ (.I(_0584_),
    .ZN(_0044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1185_ (.I(_0584_),
    .ZN(_0045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1186_ (.I(\manchester_baby_instance.BASE_0.s_tickReg ),
    .ZN(_0589_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1187_ (.A1(\manchester_baby_instance.BASE_1.s_counterValue ),
    .A2(_0589_),
    .ZN(_0590_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1188_ (.A1(\manchester_baby_instance.BASE_1.s_derivedClock ),
    .A2(_0590_),
    .Z(_0591_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1189_ (.I(_0591_),
    .Z(_0095_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1190_ (.I(_0584_),
    .ZN(_0046_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1191_ (.I(_0584_),
    .ZN(_0047_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1192_ (.I(_0584_),
    .ZN(_0048_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1193_ (.I(_0584_),
    .ZN(_0049_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1194_ (.A1(\manchester_baby_instance.BASE_1.s_counterValue ),
    .A2(_0589_),
    .Z(_0592_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1195_ (.I(_0592_),
    .Z(_0097_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1196_ (.I(\manchester_baby_instance.BASE_0.s_countReg[0] ),
    .ZN(_0098_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1197_ (.A1(_0098_),
    .A2(\manchester_baby_instance.BASE_0.s_countReg[1] ),
    .Z(_0593_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1198_ (.I(_0593_),
    .Z(_0099_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1199_ (.A1(\manchester_baby_instance.BASE_0.s_countReg[0] ),
    .A2(\manchester_baby_instance.BASE_0.s_countReg[1] ),
    .B(\manchester_baby_instance.BASE_0.s_countReg[2] ),
    .ZN(_0594_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1200_ (.I(_0594_),
    .ZN(_0100_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1201_ (.D(net74),
    .CLK(clknet_2_0__leaf_clock),
    .Q(net34),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1202_ (.D(_0000_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1203_ (.D(_0050_),
    .RN(_0001_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1204_ (.D(_0051_),
    .RN(_0002_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _1205_ (.D(_0052_),
    .RN(_0003_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _1206_ (.D(_0053_),
    .RN(_0004_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1207_ (.D(_0054_),
    .RN(_0005_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1208_ (.D(_0055_),
    .RN(_0006_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net40),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1209_ (.D(_0056_),
    .RN(_0007_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net51),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1210_ (.D(_0057_),
    .RN(_0008_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net62),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1211_ (.D(_0058_),
    .RN(_0009_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net65),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1212_ (.D(_0059_),
    .RN(_0010_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net66),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1213_ (.D(_0060_),
    .RN(_0011_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(net67),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1214_ (.D(_0061_),
    .RN(_0012_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net68),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _1215_ (.D(_0062_),
    .RN(_0013_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net69),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1216_ (.D(_0063_),
    .RN(_0014_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net70),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1217_ (.D(_0064_),
    .RN(_0015_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(net71),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1218_ (.D(_0065_),
    .RN(_0016_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(net41),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1219_ (.D(_0066_),
    .RN(_0017_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(net42),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1220_ (.D(_0067_),
    .RN(_0018_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1221_ (.D(_0068_),
    .RN(_0019_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1222_ (.D(_0069_),
    .RN(_0020_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net45),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _1223_ (.D(_0070_),
    .RN(_0021_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net46),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1224_ (.D(_0071_),
    .RN(_0022_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net47),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1225_ (.D(_0072_),
    .RN(_0023_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net48),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1226_ (.D(_0073_),
    .RN(_0024_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net49),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1227_ (.D(_0074_),
    .RN(_0025_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net50),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1228_ (.D(_0075_),
    .RN(_0026_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net52),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1229_ (.D(_0076_),
    .RN(_0027_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net53),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1230_ (.D(_0077_),
    .RN(_0028_),
    .CLK(clknet_2_1__leaf_clock),
    .Q(net54),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1231_ (.D(_0078_),
    .RN(_0029_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net55),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1232_ (.D(_0079_),
    .RN(_0030_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net56),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1233_ (.D(_0080_),
    .RN(_0031_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net57),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1234_ (.D(_0081_),
    .RN(_0032_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net58),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1235_ (.D(_0082_),
    .RN(_0033_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net59),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1236_ (.D(_0083_),
    .RN(_0034_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net60),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1237_ (.D(_0084_),
    .RN(_0035_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net61),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1238_ (.D(_0085_),
    .RN(_0036_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net63),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _1239_ (.D(_0086_),
    .RN(_0037_),
    .CLK(clknet_2_3__leaf_clock),
    .Q(net64),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1240_ (.D(_0087_),
    .RN(_0038_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1241_ (.D(_0088_),
    .RN(_0039_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1242_ (.D(_0089_),
    .RN(_0040_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1243_ (.D(_0090_),
    .RN(_0041_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1244_ (.D(_0091_),
    .RN(_0042_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _1245_ (.D(_0092_),
    .RN(_0043_),
    .CLK(clknet_2_2__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _1246_ (.D(_0093_),
    .RN(_0044_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1247_ (.D(_0094_),
    .RN(_0045_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1248_ (.D(_0095_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\manchester_baby_instance.BASE_1.s_derivedClock ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _1249_ (.D(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ),
    .RN(_0046_),
    .CLK(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ),
    .Q(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 _1250_ (.D(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[1] ),
    .RN(_0047_),
    .CLK(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ),
    .Q(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 _1251_ (.D(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[2] ),
    .RN(_0048_),
    .CLK(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ),
    .Q(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1252_ (.D(_0096_),
    .RN(_0049_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(net73),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1253_ (.D(\manchester_baby_instance.BASE_1.s_derivedClock ),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\manchester_baby_instance.BASE_1.s_bufferRegs[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1254_ (.D(_0097_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\manchester_baby_instance.BASE_1.s_counterValue ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1255_ (.D(_0098_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1256_ (.D(_0099_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1257_ (.D(_0100_),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1258_ (.D(\manchester_baby_instance.BASE_0.s_tickNext ),
    .CLK(clknet_2_0__leaf_clock),
    .Q(\manchester_baby_instance.BASE_0.s_tickReg ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clock (.I(clock),
    .Z(clknet_0_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_0__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_1__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_2__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_3__leaf_clock),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold1 (.I(\manchester_baby_instance.BASE_1.s_bufferRegs[0] ),
    .Z(net74),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1 (.I(ram_data_i[0]),
    .Z(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input10 (.I(ram_data_i[18]),
    .Z(net10),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(ram_data_i[19]),
    .Z(net11),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input12 (.I(ram_data_i[1]),
    .Z(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input13 (.I(ram_data_i[20]),
    .Z(net13),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input14 (.I(ram_data_i[21]),
    .Z(net14),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input15 (.I(ram_data_i[22]),
    .Z(net15),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input16 (.I(ram_data_i[23]),
    .Z(net16),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input17 (.I(ram_data_i[24]),
    .Z(net17),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input18 (.I(ram_data_i[25]),
    .Z(net18),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(ram_data_i[26]),
    .Z(net19),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input2 (.I(ram_data_i[10]),
    .Z(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input20 (.I(ram_data_i[27]),
    .Z(net20),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input21 (.I(ram_data_i[28]),
    .Z(net21),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input22 (.I(ram_data_i[29]),
    .Z(net22),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(ram_data_i[2]),
    .Z(net23),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input24 (.I(ram_data_i[30]),
    .Z(net24),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(ram_data_i[31]),
    .Z(net25),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(ram_data_i[3]),
    .Z(net26),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input27 (.I(ram_data_i[4]),
    .Z(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input28 (.I(ram_data_i[5]),
    .Z(net28),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input29 (.I(ram_data_i[6]),
    .Z(net29),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input3 (.I(ram_data_i[11]),
    .Z(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(ram_data_i[7]),
    .Z(net30),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input31 (.I(ram_data_i[8]),
    .Z(net31),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input32 (.I(ram_data_i[9]),
    .Z(net32),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(reset_i),
    .Z(net33),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input4 (.I(ram_data_i[12]),
    .Z(net4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input5 (.I(ram_data_i[13]),
    .Z(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(ram_data_i[14]),
    .Z(net6),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input7 (.I(ram_data_i[15]),
    .Z(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(ram_data_i[16]),
    .Z(net8),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(ram_data_i[17]),
    .Z(net9),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output34 (.I(net34),
    .Z(logisim_clock_tree_0_out),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output35 (.I(net35),
    .Z(ram_addr_o[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output36 (.I(net36),
    .Z(ram_addr_o[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(ram_addr_o[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output38 (.I(net38),
    .Z(ram_addr_o[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output39 (.I(net39),
    .Z(ram_addr_o[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output40 (.I(net40),
    .Z(ram_data_o[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output41 (.I(net41),
    .Z(ram_data_o[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output42 (.I(net42),
    .Z(ram_data_o[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output43 (.I(net43),
    .Z(ram_data_o[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output44 (.I(net44),
    .Z(ram_data_o[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output45 (.I(net45),
    .Z(ram_data_o[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output46 (.I(net46),
    .Z(ram_data_o[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output47 (.I(net47),
    .Z(ram_data_o[16]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output48 (.I(net48),
    .Z(ram_data_o[17]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output49 (.I(net49),
    .Z(ram_data_o[18]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output50 (.I(net50),
    .Z(ram_data_o[19]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output51 (.I(net51),
    .Z(ram_data_o[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output52 (.I(net52),
    .Z(ram_data_o[20]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output53 (.I(net53),
    .Z(ram_data_o[21]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output54 (.I(net54),
    .Z(ram_data_o[22]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output55 (.I(net55),
    .Z(ram_data_o[23]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output56 (.I(net56),
    .Z(ram_data_o[24]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output57 (.I(net57),
    .Z(ram_data_o[25]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output58 (.I(net58),
    .Z(ram_data_o[26]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output59 (.I(net59),
    .Z(ram_data_o[27]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output60 (.I(net60),
    .Z(ram_data_o[28]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output61 (.I(net61),
    .Z(ram_data_o[29]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output62 (.I(net62),
    .Z(ram_data_o[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output63 (.I(net63),
    .Z(ram_data_o[30]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output64 (.I(net64),
    .Z(ram_data_o[31]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output65 (.I(net65),
    .Z(ram_data_o[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output66 (.I(net66),
    .Z(ram_data_o[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output67 (.I(net67),
    .Z(ram_data_o[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output68 (.I(net68),
    .Z(ram_data_o[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output69 (.I(net69),
    .Z(ram_data_o[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output70 (.I(net70),
    .Z(ram_data_o[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output71 (.I(net71),
    .Z(ram_data_o[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output72 (.I(net72),
    .Z(ram_rw_en_o),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output73 (.I(net73),
    .Z(stop_lamp_o),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
endmodule
