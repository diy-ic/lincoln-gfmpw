module mos6502_decoder (
`ifdef USE_POWER_PINS
    inout vdd,		// User area 5.0V supply
    inout vss,		// User area ground
`endif
    input [7:0] instruction_i,
    output [65:0] decoded_instruction_o
);

    logisimTopLevelShell decoder (
        .instruction_bus_0(instruction_i[0]),
        .instruction_bus_1(instruction_i[1]),
        .instruction_bus_2(instruction_i[2]),
        .instruction_bus_3(instruction_i[3]),
        .instruction_bus_4(instruction_i[4]),
        .instruction_bus_5(instruction_i[5]),
        .instruction_bus_6(instruction_i[6]),
        .instruction_bus_7(instruction_i[7]),

        .ADC_0(decoded_instruction_o[0]),
        .AND_0(decoded_instruction_o[1]),
        .ASL_0(decoded_instruction_o[2]),
        .BCC_0(decoded_instruction_o[4]),
        .BCS_0(decoded_instruction_o[5]),
        .BEQ_0(decoded_instruction_o[6]),
        .BMI_0(decoded_instruction_o[7]),
        .BNE_0(decoded_instruction_o[8]),
        .BPL_0(decoded_instruction_o[9]),
        .BRK_0(decoded_instruction_o[10]),
        .BVC_0(decoded_instruction_o[11]),
        .BVS_0(decoded_instruction_o[12]),
        .CLC_0(decoded_instruction_o[13]),
        .CLD_0(decoded_instruction_o[14]),
        .CLI_0(decoded_instruction_o[15]),
        .CLV_0(decoded_instruction_o[16]),
        .CMP_0(decoded_instruction_o[17]),
        .CPX_0(decoded_instruction_o[18]),
        .CPY_0(decoded_instruction_o[19]),
        .DEC_0(decoded_instruction_o[20]),
        .DES_0(decoded_instruction_o[21]),
        .DEY_0(decoded_instruction_o[22]),
        .EOR_0(decoded_instruction_o[23]),
        .INC_0(decoded_instruction_o[24]),
        .INX_0(decoded_instruction_o[25]),
        .INY_0(decoded_instruction_o[26]),
        .JMP_0(decoded_instruction_o[27]),
        .JSR_0(decoded_instruction_o[28]),
        .LDA_0(decoded_instruction_o[29]),
        .LDX_0(decoded_instruction_o[30]),
        .LDX_Y_0(decoded_instruction_o[31]),
        .LDY_0(decoded_instruction_o[32]),
        .LSR_0(decoded_instruction_o[33]),
        .ORA_0(decoded_instruction_o[34]),
        .PHA_0(decoded_instruction_o[35]),
        .PHP_0(decoded_instruction_o[36]),
        .PLA_0(decoded_instruction_o[37]),
        .PLP_0(decoded_instruction_o[38]),
        .ROL_0(decoded_instruction_o[39]),
        .ROR_0(decoded_instruction_o[40]),
        .RTI_0(decoded_instruction_o[41]),
        .RTS_0(decoded_instruction_o[42]),
        .SBC_0(decoded_instruction_o[43]),
        .SEC_0(decoded_instruction_o[44]),
        .SED_0(decoded_instruction_o[45]),
        .SEI_0(decoded_instruction_o[46]),
        .STA_0(decoded_instruction_o[47]),
        .STX_0(decoded_instruction_o[48]),
        .STY_0(decoded_instruction_o[49]),
        .TAX_0(decoded_instruction_o[50]),
        .TAY_0(decoded_instruction_o[51]),
        .TKA_0(decoded_instruction_o[52]),
        .TKS_0(decoded_instruction_o[53]),
        .TSX_0(decoded_instruction_o[54]),
        .TYA_0(decoded_instruction_o[55]),
        .A_0(decoded_instruction_o[3]),
        .Xind_0(decoded_instruction_o[56]),
        .absX_0(decoded_instruction_o[57]),
        .absY_0(decoded_instruction_o[58]),
        .abs_0(decoded_instruction_o[59]),
        .hash_0(decoded_instruction_o[60]),
        .indY_0(decoded_instruction_o[61]),
        .ind_0(decoded_instruction_o[62]),
        .rel_0(decoded_instruction_o[63]),
        .zpgX_0(decoded_instruction_o[64]),
        .zpg_0(decoded_instruction_o[65])
    );

endmodule